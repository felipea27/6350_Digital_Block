##################################################################################
#
#           GLOBALFOUNDRIES
#
#     22FDSOI EDI/Innovus technology file
#
##################################################################################

####################################################################################
#
# ----------------------------- DISCLAIMER -----------------------------------------
# EDI Version - complete Innovus behavior not analyzed yet !    
#
####################################################################################

#==============================================================================
# Revision: 1.0_2.5
# Date: 23 January 2025
#-------------------------------------------------------
# target: 22FDSOI process
# metal stack: 10M_2Mx_5Cx_1Jx_2Qx_LB
# site: unit must be defined in std-cell.lef
# first vertical pitch based on Critical-Poly-Pitch: 116cpp
# editor: GF 
# Preferred routing directions:
# vertical:   M1 C1 C3 C5 QA LB 
# horizontal: M2 C2 C4 JA QB
#------------------------------------------------------
# Known Issues
# - inter-VT spacing is not enabled due to missing support of allowed abutment
# - property EDGETYPE is defined just to support related reference library constraints 
# - Cx T2T extension pessimism (23 -> 46nm) is due to Innovus 15.12.00 behavior (GF-Bug-030773)
# - we do not limit the via number to 128 as long as no urgent via got automatically removed (S-Router-WARNING)
# - combination of PARALLELRUNLENGTH spacing table and TWOWIDTHS spacing table for Mx with minor pessimism
# - no support of special new 30x/34x PAD rules
# - warnings regarding minWidth violations in JQ vias can be ignored
# - 7.5t variant of STD-Libs need special track definitions (B-236952) during floorplanning:
#    add_tracks -pitch_pattern {{M2 offset 0.06 {pitch 0.08 repeat 6} pitch 0.12}} 
# - no support of minArea rules for fill shapes if those are on standard metal (MxEz.A.3 vs. CFOMxEz.A.1 ) - see B-262387
# - if customer need to use tool version older than 19.13 - you need to switch CB TYPE back to MASTERSLICE 
# - modified Mx OFFSET depending on used std-cell library may help to to get better pin access or 100% multi cut usage






#--------------------------------------------------------------------------------
# Note: Required tool version / Evaluated with Innovus 22.13.000
#--------------------------------------------------------------------------------

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;
CLEARANCEMEASURE EUCLIDEAN ;
# USEMINSPACING OBS OFF ;  Customer can change the settings due to IP/macro blockage/OBS generation style
USEMINSPACING OBS ON ;

PROPERTYDEFINITIONS
  MACRO oaTaper STRING ;
  MACRO vceLastSavedModifiedCounter INTEGER ;
  MACRO LEF58_EDGETYPE STRING ; 
    LAYER LEF58_MINSTEP STRING ;
    LAYER LEF58_SPACING STRING ;
    LAYER LEF58_AREA STRING ;
    LAYER LEF58_CUTCLASS STRING ;
    LAYER LEF58_ENCLOSURE STRING ;
    LAYER LEF58_ENCLOSURETOJOINT STRING ;
    LAYER LEF58_MINIMUMCUT STRING ;
    LAYER LEF58_MINWIDTH STRING ;
    LAYER LEF58_VIACLUSTER STRING ;
    LAYER LEF58_ARRAYSPACING STRING ;
    LAYER LEF58_SPACINGTABLE STRING ;
    LAYER LEF58_ENCLOSUREEDGE STRING ;
    LAYER LEF58_EOLEXTENSIONSPACING STRING ;
    LAYER LEF58_ENCLOSUREWIDTH STRING ;
    LAYER LEF58_WIDTHTABLE STRING ;
    LAYER LEF58_WIDTH STRING ;
    LAYER LEF58_VOLTAGESPACING STRING ;
    LAYER LEF58_EOLENCLOSURE STRING ;
    LAYER LEF57_ANTENNAGATEPLUSDIFF STRING ;
    LAYER LEF58_TYPE STRING ;
    LAYER LEF58_JOINTCORNERSPACING STRING ;
    LAYER LEF58_FORBIDDENSPACING STRING ;
    LAYER LEF58_TWOWIRESFORBIDDENSPACING STRING ;

    LIBRARY LEF58_CELLEDGESPACINGTABLE STRING
    "CELLEDGESPACINGTABLE
        EDGETYPE BOTHDRAIN BOTHDRAIN 0.348
        EDGETYPE BOTHDRAIN SOURCEDRAIN 0.348
        EDGETYPE BOTHDRAIN DRAINSOURCE 0.348
        EDGETYPE BOTHDRAIN BOTHSOURCE 0.000
        EDGETYPE BOTHSOURCE BOTHSOURCE 0.000
        EDGETYPE BOTHSOURCE DRAINSOURCE 0.000
        EDGETYPE BOTHSOURCE SOURCEDRAIN 0.000
        EDGETYPE DRAINSOURCE DRAINSOURCE 0.348
        EDGETYPE SOURCEDRAIN SOURCEDRAIN 0.348
        EDGETYPE SOURCEDRAIN DRAINSOURCE 0.000
	EDGETYPE SC8T_116CPP_BASE_CSC_SOURCE       SC8T_116CPP_BASE_CSC_SOURCE	   EXCEPTABUTTED   0.232
	EDGETYPE SC8T_116CPP_BASE_CSC_DRAIN        SC8T_116CPP_BASE_CSC_SOURCE	   EXCEPTABUTTED   0.232
	EDGETYPE SC8T_116CPP_BASE_CSC_DRAIN        SC8T_116CPP_BASE_CSC_DRAIN	                   0.116
	EDGETYPE SC8T_116CPP_BASE_CSC_SOURCE2CPP   SC8T_116CPP_BASE_CSC_SOURCE2CPP   EXCEPTABUTTED   0.232
	EDGETYPE SC8T_116CPP_BASE_CSC_SOURCE       SC8T_116CPP_BASE_CSC_SOURCE2CPP   EXCEPTABUTTED   0.232
	EDGETYPE SC8T_116CPP_BASE_CSC_SOURCE2CPP   SC8T_116CPP_BASE_CSC_DRAIN	                   0.232
	EDGETYPE SC7P5T_116CPP_BASE_CSC_SOURCE     SC7P5T_116CPP_BASE_CSC_SOURCE     EXCEPTABUTTED   0.232 
	EDGETYPE SC7P5T_116CPP_BASE_CSC_DRAIN      SC7P5T_116CPP_BASE_CSC_SOURCE     EXCEPTABUTTED   0.232 
	EDGETYPE SC7P5T_116CPP_BASE_CSC_DRAIN      SC7P5T_116CPP_BASE_CSC_DRAIN                      0.116 
	EDGETYPE SC7P5T_116CPP_BASE_CSC_SOURCE2CPP SC7P5T_116CPP_BASE_CSC_SOURCE2CPP EXCEPTABUTTED   0.232
	EDGETYPE SC7P5T_116CPP_BASE_CSC_SOURCE     SC7P5T_116CPP_BASE_CSC_SOURCE2CPP EXCEPTABUTTED   0.232
	EDGETYPE SC7P5T_116CPP_BASE_CSC_SOURCE2CPP SC7P5T_116CPP_BASE_CSC_DRAIN                      0.232
	EDGETYPE SC12T_116CPP_BASE_CSC_SOURCE       SC12T_116CPP_BASE_CSC_SOURCE     EXCEPTABUTTED   0.232
	EDGETYPE SC12T_116CPP_BASE_CSC_DRAIN        SC12T_116CPP_BASE_CSC_SOURCE     EXCEPTABUTTED   0.232
	EDGETYPE SC12T_116CPP_BASE_CSC_DRAIN        SC12T_116CPP_BASE_CSC_DRAIN                      0.116
	EDGETYPE SC12T_116CPP_BASE_CSC_SOURCE2CPP   SC12T_116CPP_BASE_CSC_SOURCE2CPP EXCEPTABUTTED   0.232
	EDGETYPE SC12T_116CPP_BASE_CSC_SOURCE       SC12T_116CPP_BASE_CSC_SOURCE2CPP EXCEPTABUTTED   0.232
	EDGETYPE SC12T_116CPP_BASE_CSC_SOURCE2CPP   SC12T_116CPP_BASE_CSC_DRAIN                      0.232
      ;" ;
 
END PROPERTYDEFINITIONS

#--------------------------------------------------------------------------------
# No Site definition in tech.lef - need to be defined in std-cell.lef
#--------------------------------------------------------------------------------


################################################# VT ############################################

LAYER LVTN
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;  
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END LVTN
LAYER LVTP
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
#  SPACING 0.208 LAYER LVTN ;  removed as workaround because abutment is alowed
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END LVTP

LAYER SLVTN
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
#  SPACING 0.208 LAYER LVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER LVTP ;  removed as workaround because abutment is alowed
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END SLVTN
LAYER SLVTP
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
#  SPACING 0.208 LAYER LVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER LVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTN ;  removed as workaround because abutment is alowed
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END SLVTP

LAYER RVTN
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
#  SPACING 0.208 LAYER LVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER LVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTP ;  removed as workaround because abutment is alowed
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END RVTN
LAYER RVTP
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
#  SPACING 0.208 LAYER LVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER LVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER RVTN ;  removed as workaround because abutment is alowed
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END RVTP

LAYER HVTN
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
#  SPACING 0.208 LAYER LVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER LVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER RVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER RVTP ;  removed as workaround because abutment is alowed
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END HVTN
LAYER HVTP
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
#  SPACING 0.208 LAYER LVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER LVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER SLVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER RVTN ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER RVTP ;  removed as workaround because abutment is alowed
#  SPACING 0.208 LAYER HVTN ;  removed as workaround because abutment is alowed
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END HVTP

LAYER LLN
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END LLN
LAYER LLP
  TYPE IMPLANT ;
  SPACING 0.208 ;
#  WIDTH 0.208 ;    
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;  
END LLP

LAYER ULLN
  TYPE IMPLANT ;
  SPACING 0.232 ;
#  WIDTH 0.232 ;    
  PROPERTY LEF58_AREA "
    AREA   0.071 ; " ;  
END ULLN
LAYER ULLP
  TYPE IMPLANT ;
  SPACING 0.232 ;
#  WIDTH 0.232 ;    
  PROPERTY LEF58_AREA "
    AREA   0.071 ; " ;  
END ULLP
LAYER EGSLVTN
  TYPE IMPLANT ;
  SPACING 0.208 ;
  PROPERTY LEF58_AREA "
    AREA   0.064 ; " ;
END EGSLVTN
LAYER EGSLVTP
  TYPE IMPLANT ;
  SPACING 0.208 ;
  PROPERTY LEF58_AREA "
    AREA   0.198 ; " ;
END EGSLVTP
LAYER EGLVTN
  TYPE IMPLANT ;
  SPACING 0.208 ;
  PROPERTY LEF58_AREA "
    AREA   0.198 ; " ;
END EGLVTN
LAYER EGLVTP
  TYPE IMPLANT ;
  SPACING 0.208 ;
  PROPERTY LEF58_AREA "
    AREA   0.198 ; " ;
END EGLVTP
LAYER EGULLP
  TYPE IMPLANT ;
  SPACING 0.208 ;
  PROPERTY LEF58_AREA "
    AREA   0.198 ; " ;
END EGULLP

LAYER EGUOSLVTN
  TYPE IMPLANT ;
  SPACING 0.208 ;
  PROPERTY LEF58_AREA "
    AREA   0.198 ; " ;
END EGUOSLVTN


LAYER LV
  TYPE MASTERSLICE ;
END LV

LAYER RS
  TYPE MASTERSLICE ;
END RS


################### Marker layer 7t and 6.75t for FDX-EXT, MK7 for FDX ##########################

LAYER CLIB_MKR1
    TYPE MASTERSLICE ;
END CLIB_MKR1 

LAYER CLIB_MKR4
    TYPE MASTERSLICE ;
END CLIB_MKR4 

LAYER CLIB_MKR41
    TYPE MASTERSLICE ;
END CLIB_MKR41 

LAYER CLIB_MKR5
    TYPE MASTERSLICE ;
END CLIB_MKR5 

LAYER CLIB_MKR51
    TYPE MASTERSLICE ;
END CLIB_MKR51 

LAYER CLIB_MKR3
    TYPE MASTERSLICE ;
END CLIB_MKR3

LAYER CLIB_MKR61
    TYPE MASTERSLICE ;
END CLIB_MKR61

LAYER MIXVT
    TYPE MASTERSLICE ;
END MIXVT

################################################# FEOL #########################################

LAYER RX
    TYPE MASTERSLICE ;
    PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
END RX

LAYER NW
    TYPE MASTERSLICE ;
    PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END NW

LAYER SXCUT
    TYPE MASTERSLICE ;
    PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END SXCUT

LAYER PC
    TYPE MASTERSLICE ;
END PC

LAYER CB
    TYPE CUT ;
END CB

LAYER CA
    TYPE CUT ;
END CA

################################################## BEOL ###########################################


LAYER M1
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION VERTICAL ;
  PITCH 0.116 0.080 ;
  OFFSET   0.058 0.000 ;
# M1Ez.W.1
    MINWIDTH 0.040 ;

# M1Ez.W.2
    MAXWIDTH 1.700 ;

# M1Ez.W.1
    WIDTH    0.040 ;

# M1Ez.A.5
    MINENCLOSEDAREA 0.160 ; 

# M1Ez.A.2
    AREA     0.0064 ;

# M1Ez.A.1
    PROPERTY LEF58_AREA "AREA 0.0074 EXCEPTRECTANGLE ; " ;

# M1Ez.SE.1   ?? SE.2
    MINSTEP 0.057 MAXEDGES 1 ; 

# MxEz.SE.2
    PROPERTY LEF58_MINSTEP "
       MINSTEP 0.02 MAXEDGES 1 MINADJACENTLENGTH 0.07 ; " ;

# M1Ez.S.1
    PROPERTY LEF58_SPACING "SPACING 0.060 SAMEMASK ; " ;

# M1Ez.S.3 diff mask
    SPACING 0.040 ;

# M1Ez.S.3/14/17 diff mask
  SPACINGTABLE  TWOWIDTHS
			   ###     width=  0.000  0.072  0.120   0.156   0.208 
			   ###     prl=    none   0.000  0.000   0.000   0.300 
			   ###     ---------------------------------------------
		WIDTH 0.000                0.040  0.040  0.050   0.054   0.090 
		WIDTH 0.072 PRL 0.000      0.040  0.040  0.050   0.054   0.090 
		WIDTH 0.120 PRL 0.000      0.050  0.050  0.050   0.054   0.090 
		WIDTH 0.156 PRL 0.000      0.054  0.054  0.054   0.054   0.090 
		WIDTH 0.208 PRL 0.300      0.090  0.090  0.090   0.090   0.090  ;


# first part: M1Ez.S.1/8/9/14-20 same mask - Pessimistic support for M1Ez.S.8/9 due to PRL increase condition
# second part: M1Ez.S.1/1a/2/8/9/10/14-20 same mask --> removed due to WARNING (NRDB-947)
  PROPERTY LEF58_SPACINGTABLE  "
  SPACINGTABLE  TWOWIDTHS  SAMEMASK
		WIDTH 0.000                0.060   0.060   0.066   0.066  0.100  0.100 
		WIDTH 0.072 PRL 0.000      0.060   0.060   0.066   0.074  0.100  0.103 
		WIDTH 0.080 PRL 0.080      0.066   0.066   0.066   0.074  0.100  0.103 
		WIDTH 0.156 PRL 0.000      0.066   0.074   0.074   0.082  0.100  0.111 
		WIDTH 0.159 PRL 0.160      0.100   0.100   0.100   0.100  0.100  0.111 
		WIDTH 0.208 PRL 0.300      0.100   0.103   0.103   0.111  0.111  0.140  ; " ; 

# M1Ez.S.4/5 same mask T2L and T2T
    PROPERTY LEF58_SPACING "
        SPACING 0.070 ENDOFLINE 0.060 WITHIN 0.020 SAMEMASK ENDTOEND 0.080 EXTENSION 0.020 MINLENGTH 0.001 TWOSIDES ; " ;

# M1Ez.S.5/6: diff mask  T2L and T2T
    PROPERTY LEF58_SPACING "
        SPACING 0.040 ENDOFLINE 0.060 WITHIN 0.020 ENDTOEND 0.040 EXTENSION 0.020 MINLENGTH 0.001 TWOSIDES ; " ;

# M1Ez.S.19
#    PROPERTY LEF58_SPACING "
#        SPACING 0.065 ENDOFLINE 0.046 OPPOSITEWIDTH 0.038 WITHIN 0.009 SAMEMASK ENDTOEND 0.08 MINLENGTH 0.020 TWOSIDES ; " ;
# M1Ez.S.21
# this rule says width <= 0.038
#   PROPERTY LEF58_SPACING "
#       SPACING 0.075 ENDOFLINE 0.039 OPPOSITEWIDTH 0.048 WITHIN 0.016 PARALLELEDGE 0.066 WITHIN 0.050 TWOEDGES ; " ;  


# Vx.C.15 # Vx.C.12/13/14
    PROPERTY LEF58_MINIMUMCUT "
        MINIMUMCUT CUTCLASS Vx 2  WIDTH 0.185 WITHIN 0.221 FROMABOVE ;
        MINIMUMCUT CUTCLASS Vx 3  WIDTH 0.349 WITHIN 0.221 FROMABOVE ;
        MINIMUMCUT CUTCLASS Vx 4  WIDTH 0.479 WITHIN 0.221 FROMABOVE ;
        MINIMUMCUT  CUTCLASS VxBAR 1 WIDTH 0.185 WITHIN 0.181 FROMABOVE ;
        MINIMUMCUT  CUTCLASS VxBAR 2 WIDTH 0.349 WITHIN 0.181 FROMABOVE ;
        MINIMUMCUT  CUTCLASS VxBAR 2 WIDTH 0.479 WITHIN 0.181 FROMABOVE ;
        MINIMUMCUT CUTCLASS Vx 2 WIDTH 0.185 WITHIN 0.221 FROMABOVE LENGTH 0.186 WITHIN 1.401 ; " ;



# M1Ez.S.32-41
    PROPERTY LEF58_VOLTAGESPACING
     "VOLTAGESPACING
     1.32 0.045
     1.65 0.050
     1.98 0.060
     2.75 0.070
     3.63 0.100 
     5.50 0.120
     7.70 0.150
     11.0 0.180
     16.5 0.200
     18.7 0.220 ; " ;


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END M1


LAYER V1
  TYPE CUT ;

# Vx.LW.1 # VxBAR.W.1, VxBAR.L.1 
    PROPERTY LEF58_CUTCLASS "
        CUTCLASS Vx    WIDTH 0.040              CUTS 1 ;
        CUTCLASS VxBAR WIDTH 0.040 LENGTH 0.080 CUTS 2 ; " ;

# Vx.C.1 SAVx
  PROPERTY LEF58_ENCLOSUREEDGE "
    ENCLOSUREEDGE CUTCLASS Vx ABOVE 0.005 OPPOSITE ; " ;
# Vx.C.3/4 SAVx
  PROPERTY LEF58_VIACLUSTER "
    VIACLUSTER CUTCLASS Vx CUTS 0 DIAGONAL 5 WITHIN 0.040 0.046 ; " ;

# Vx.S.3,  Vx.S.1d,      Vx.S.VxBAR2, Vx.S.VxBAR.1, VxLRG.S.Vx.1 
# Vx.S.VxBAR.2, VxBAR.S.1a/2a, VxLRG.S.VxBAR.1
# Vx.S.VxBAR.1, VxBAR.S.2a, VxBAR.S.1b,  VxLRG.S.VxBAR.2
# VxBAR.S.1b = 0.072 with extension of 0.020. However we are going with the conservation value of 0.112 since we dont have syntax for it.

    PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
        CENTERANDEDGE  Vx TO Vx
        CUTCLASS          Vx        VxBAR SIDE     VxBAR END
        Vx          0.113  0.075  0.072  0.090  0.072  0.090
        VxBAR SIDE  0.072  0.090  0.080  0.080  0.100  0.100
        VxBAR END   0.072  0.090  0.100  0.100  0.100  0.100 ; " ;

# Vx.C.5 The maximum number of neighboring Vx at center to center space <0.130um, z=1-2.  <=2 
  PROPERTY LEF58_SPACING "
    SPACING 0.130 CENTERTOCENTER ADJACENTCUTS 3 WITHIN 0.130 CUTCLASS Vx ; " ;

#Vx.EX.MxEz.1.or.a/b/c, Vx.EX.MyEz.1.or.a/b/c 
#Vx.Ex.MxEz.2, Vx.EZ.MyEz.2
#Vx.EN.MyEz.2
#Vx.EX.MxEz.4.or.a, Vx.EN.MyEz.3
#Vx.EN.MyEz.4
#Vx.EN.MxEz.5, Vx.EN.MyEz.5
#Vx.EN.MxEz.6
#Vx.EN.MxEz.7, Vx.EN.MyEz.7
#VxBAR.EX.MxEz.1.or.a/b/c, VxBAR.EX.MyEz.1.or.a/b/c
#VxBAR.EN.MxEz.3, VxBAR.EN.MyEz.2
#VxBAR.EN.MxEz.4, VxBAR.EN.MyEz.3
#VxBAR.EN.MyEz.4
#VxBAR.EN.MxEz.5, VxBAR.EN.MyEz.5
#VxBAR.EN.MxEz.6
#VxBAR.EN.MxEz.7, VxBAR.EN.MyEz.7
#
    PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS Vx       0.000 0.030 ;
    ENCLOSURE CUTCLASS Vx       0.007 0.025 ;
    ENCLOSURE CUTCLASS Vx BELOW 0.010 0.020 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.020 0.020 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.003 0.030 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.007 0.025 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.020 0.020 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.005 0.030 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.007 0.025 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.020 0.020 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.010 0.025 WIDTH 0.060 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.020 0.020 WIDTH 0.060 ;
    ENCLOSURE CUTCLASS Vx BELOW 0.010 0.020 WIDTH 0.080 ;
    ENCLOSURE CUTCLASS Vx ABOVE 0.020 0.020 WIDTH 0.080 ;
    ENCLOSURE CUTCLASS Vx BELOW 0.020 0.020 WIDTH 0.120 ;
    ENCLOSURE CUTCLASS Vx       0.025 0.025 WIDTH 0.200 ;
    ENCLOSURE CUTCLASS VxBAR END 0.000 SIDE 0.030 ;
    ENCLOSURE CUTCLASS VxBAR END 0.030 SIDE 0.000 ;
    ENCLOSURE CUTCLASS VxBAR END 0.007 SIDE 0.025 ;
    ENCLOSURE CUTCLASS VxBAR END 0.025 SIDE 0.007 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.010 SIDE 0.020 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.020 SIDE 0.010 ;
    ENCLOSURE CUTCLASS VxBAR ABOVE END 0.020 SIDE 0.020 ;
    ENCLOSURE CUTCLASS VxBAR END 0.003 SIDE 0.030 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS VxBAR END 0.030 SIDE 0.003 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS VxBAR END 0.007 SIDE 0.025 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS VxBAR END 0.025 SIDE 0.007 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS VxBAR ABOVE END 0.020 SIDE 0.020 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.010 SIDE 0.020 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.020 SIDE 0.010 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS VxBAR END 0.005 SIDE 0.030 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VxBAR END 0.030 SIDE 0.005 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VxBAR END 0.007 SIDE 0.025 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VxBAR END 0.025 SIDE 0.007 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VxBAR ABOVE END 0.020 SIDE 0.020 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.010 SIDE 0.020 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.020 SIDE 0.010 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VxBAR ABOVE END 0.010 SIDE 0.025 WIDTH 0.060 ;
    ENCLOSURE CUTCLASS VxBAR ABOVE END 0.025 SIDE 0.010 WIDTH 0.060 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.010 SIDE 0.020 WIDTH 0.080 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.020 SIDE 0.010 WIDTH 0.080 ;
    ENCLOSURE CUTCLASS VxBAR ABOVE END 0.020 SIDE 0.020 WIDTH 0.080 ;
    ENCLOSURE CUTCLASS VxBAR BELOW END 0.020 SIDE 0.020 WIDTH 0.120 ;
    ENCLOSURE CUTCLASS VxBAR END 0.030 SIDE 0.030 WIDTH 0.200 ;
    ENCLOSURE CUTCLASS VxBAR END 0.030 SIDE 0.030 WIDTH 0.200 ; " ;
		
# Vx.EX.MxEz/MyEz.2
    PROPERTY LEF58_EOLENCLOSURE "
    EOLENCLOSURE 0.105 CUTCLASS Vx BELOW 0.010 MINLENGTH 0.021 ;
    EOLENCLOSURE 0.105 CUTCLASS Vx ABOVE 0.020 MINLENGTH 0.021 ; " ;
		
# Vx.S.MyEz.1, VxBAR.S.MyEz.1
  PROPERTY LEF58_SPACING "
	SPACING 0.02 LAYER M2 CUTCLASS Vx CONCAVECORNER ; " ;
  PROPERTY LEF58_SPACING "
	SPACING 0.02 LAYER M2 CUTCLASS VxBAR CONCAVECORNER ; " ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END V1


LAYER M2 
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.080 0.080 ;
  OFFSET    0.080 0.080 ;

# MxEz.W.1
    MINWIDTH 0.040 ;

# MxEz.W.2
    MAXWIDTH 1.700 ;

# MxEz.W.1
    WIDTH    0.040 ;

# MxEz.A.5
    MINENCLOSEDAREA 0.160 ; 

# MxEz.A.2
    AREA     0.0088 ;

# MxEz.A.1
    PROPERTY LEF58_AREA "AREA 0.011 EXCEPTRECTANGLE ; " ;

# MxEz.A.3 greater/equal 0.060
PROPERTY LEF58_AREA
       "AREA 0.0088 RECTWIDTH 0.059 ;
        AREA 0.0110 RECTWIDTH 1.700 ; " ;

# MxEz.SE.1   ?? SE.2
    MINSTEP 0.057 MAXEDGES 1 ; 
    
# MxEz.SE.2
    PROPERTY LEF58_MINSTEP "
       MINSTEP 0.02 MAXEDGES 1 MINADJACENTLENGTH 0.08 ; " ;

# MxEz.S.1
    PROPERTY LEF58_SPACING "SPACING 0.060 SAMEMASK ; " ;

# MxEz.S.3 diff mask
    SPACING 0.040 ;

# MxEz.S.12 
    PROPERTY LEF58_SPACING "
       SPACING 0.080 NOTCHLENGTH 0.120 NOTCHWIDTH 0.049 ; " ;

# MxEz.S.3a
    SPACING 0.064 NOTCHLENGTH 0.000 ;

 # MxEz.S.3/13-20 diff mask
  SPACINGTABLE  TWOWIDTHS
			   ###     width=  0.000  0.072  0.120   0.156   0.208 
			   ###     prl=    none   0.000  0.000   0.000   0.300 
			   ###     ---------------------------------------------
		WIDTH 0.000                0.040  0.040  0.050   0.066   0.090 
		WIDTH 0.072 PRL 0.000      0.040  0.040  0.050   0.074   0.090 
		WIDTH 0.120 PRL 0.000      0.050  0.050  0.050   0.074   0.090 
		WIDTH 0.156 PRL 0.000      0.066  0.074  0.074   0.082   0.090 
		WIDTH 0.208 PRL 0.300      0.090  0.090  0.090   0.090   0.090  ;


# MxEz.S.1/1a/2/8/9/10/14-20 same mask 
  PROPERTY LEF58_SPACINGTABLE  "
  SPACINGTABLE  TWOWIDTHS  SAMEMASK
		WIDTH 0.000                0.060  0.064  0.080 0.060  0.068  0.068 0.068  0.100  0.100 
		WIDTH 0.000 PRL 0.700      0.064  0.064  0.080 0.064  0.068  0.068 0.074  0.100  0.100 
		WIDTH 0.000 PRL 2.999      0.080  0.080  0.080 0.080  0.080  0.080 0.080  0.100  0.100 
		WIDTH 0.072 PRL 0.000      0.060  0.064  0.080 0.060  0.068  0.068 0.074  0.100  0.103 
		WIDTH 0.080 PRL 0.000      0.068  0.068  0.080 0.068  0.068  0.068 0.074  0.100  0.103 
		WIDTH 0.099 PRL 0.000      0.068  0.068  0.080 0.068  0.068  0.080 0.080  0.100  0.103 
		WIDTH 0.156 PRL 0.000      0.068  0.068  0.080 0.074  0.074  0.080 0.082  0.100  0.111 
		WIDTH 0.159 PRL 0.160      0.100  0.100  0.100 0.100  0.100  0.100 0.100  0.100  0.111 
		WIDTH 0.208 PRL 0.300      0.100  0.100  0.100 0.103  0.103  0.103 0.111  0.111  0.140  ; " ;

# MxEz.S.11 corner spacing - same mask		       
  PROPERTY LEF58_JOINTCORNERSPACING "
    JOINTCORNERSPACING 0.077 SAMEMASK JOINTWIDTH 0.080 MINLENGTH 0.02 JOINTLENGTH 0.056 EDGELENGTH 0.056 ; " ;

# MxEz.S.4/5 same mask T2L and T2T
    PROPERTY LEF58_SPACING "
        SPACING 0.070 ENDOFLINE 0.060 WITHIN 0.020 SAMEMASK ENDTOEND 0.080 EXTENSION 0.020 MINLENGTH 0.001 TWOSIDES ; " ;

# MxEz.S.5/6: diff mask  T2L and T2T
    PROPERTY LEF58_SPACING "
        SPACING 0.040 ENDOFLINE 0.060 WITHIN 0.020 ENDTOEND 0.040 EXTENSION 0.020 MINLENGTH 0.001 TWOSIDES ; " ;


# AY/Vx.C.12/13/14/15
    PROPERTY LEF58_MINIMUMCUT "
        MINIMUMCUT CUTCLASS Vx 2  WIDTH 0.185 WITHIN 0.221 FROMBELOW  ;
        MINIMUMCUT CUTCLASS Vx 3  WIDTH 0.349 WITHIN 0.221 FROMBELOW  ;
        MINIMUMCUT CUTCLASS Vx 4  WIDTH 0.479 WITHIN 0.221 FROMBELOW  ;
        MINIMUMCUT  CUTCLASS VxBAR 1 WIDTH 0.185 WITHIN 0.181 FROMBELOW  ;
        MINIMUMCUT  CUTCLASS VxBAR 2 WIDTH 0.349 WITHIN 0.181 FROMBELOW  ;
        MINIMUMCUT  CUTCLASS VxBAR 2 WIDTH 0.479 WITHIN 0.181 FROMBELOW  ;
        MINIMUMCUT CUTCLASS Vx 2 WIDTH 0.185 WITHIN 0.221 FROMBELOW  LENGTH 0.186 WITHIN 1.401 ;  
        MINIMUMCUT CUTCLASS AY 2  WIDTH 0.185 WITHIN 0.221  FROMABOVE ;
        MINIMUMCUT CUTCLASS AY 3  WIDTH 0.349 WITHIN 0.221 FROMABOVE ;
        MINIMUMCUT CUTCLASS AY 4  WIDTH 0.479 WITHIN 0.221 FROMABOVE ;
        MINIMUMCUT  CUTCLASS AYBAR 1 WIDTH 0.185 WITHIN 0.181  FROMABOVE ;
        MINIMUMCUT  CUTCLASS AYBAR 2 WIDTH 0.349 WITHIN 0.181  FROMABOVE ;
        MINIMUMCUT  CUTCLASS AYBAR 2 WIDTH 0.479 WITHIN 0.181  FROMABOVE ;
        MINIMUMCUT CUTCLASS AY 2 WIDTH 0.185 WITHIN 0.221 FROMABOVE LENGTH 0.186 WITHIN 1.401 ; " ;  



# MxEz.S.32-41
    PROPERTY LEF58_VOLTAGESPACING
     "VOLTAGESPACING
     1.32 0.045
     1.65 0.050
     1.98 0.060
     2.75 0.070
     3.63 0.100 
     5.50 0.120
     7.70 0.150
     11.0 0.180
     16.5 0.200
     18.7 0.220 ; " ;


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END M2

LAYER AY
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
    CUTCLASS AY    WIDTH 0.040 ;
    CUTCLASS AYBAR WIDTH 0.040 LENGTH 0.080 CUTS 2 ; " ;

# AY.S... - AY minimum space to AY for runlength > 0 um and < 0.040um 
  PROPERTY LEF58_SPACINGTABLE "
     SPACINGTABLE
       CENTERANDEDGE AY TO AY
        CUTCLASS          AY        AYBAR SIDE     AYBAR END       
         AY         0.120  0.090  0.072  0.090  0.072  0.090 
        AYBAR SIDE  0.072  0.090  0.080  0.080  0.100  0.100 
        AYBAR END   0.072  0.090  0.100  0.100  0.100  0.100 ; " ;

# AY.C.1 The mAYimum number of neighboring AY at center to center space <0.127um, z=1-2.  <=2 
  PROPERTY LEF58_SPACING "
    SPACING 0.127 CENTERTOCENTER ADJACENTCUTS 3 WITHIN 0.127 CUTCLASS AY ; " ;

# AY.EN....
  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS AY BELOW 0.000 0.030 ;
    ENCLOSURE CUTCLASS AY BELOW 0.007 0.025 ;
    ENCLOSURE CUTCLASS AY       0.020 0.020 ;
    ENCLOSURE CUTCLASS AY ABOVE 0.002 0.034 ; 
    ENCLOSURE CUTCLASS AY ABOVE 0.007 0.030 ; 
    ENCLOSURE CUTCLASS AY	0.030 0.030 WIDTH 0.200 ;
    ENCLOSURE CUTCLASS AY BELOW 0.020 0.020 WIDTH 0.100 ; 
    ENCLOSURE CUTCLASS AY BELOW 0.010 0.025 WIDTH 0.080 ; 
    ENCLOSURE CUTCLASS AY BELOW 0.020 0.020 WIDTH 0.080 ; 
    ENCLOSURE CUTCLASS AY BELOW 0.005 0.030 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS AY BELOW 0.007 0.025 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS AY BELOW 0.003 0.030 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS AY BELOW 0.007 0.025 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS AY ABOVE 0.005 0.034 WIDTH 0.051 ; 
    ENCLOSURE CUTCLASS AY ABOVE 0.007 0.030 WIDTH 0.051 ;	  
    ENCLOSURE CUTCLASS AY ABOVE 0.020 0.020 WIDTH 0.051 ; 
    ENCLOSURE CUTCLASS AY ABOVE 0.010 0.030 WIDTH 0.060 ;	  
    ENCLOSURE CUTCLASS AY ABOVE 0.020 0.020 WIDTH 0.060 ; 
    ENCLOSURE CUTCLASS AY ABOVE 0.020 0.020 WIDTH 0.080 ;	  
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.000 SIDE 0.030 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.030 SIDE 0.000 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.007 SIDE 0.025 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.025 SIDE 0.007 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.010 SIDE 0.020 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.020 SIDE 0.010 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.003 SIDE 0.030 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.030 SIDE 0.003 WIDTH 0.046 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.005 SIDE 0.030 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.030 SIDE 0.005 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.010 SIDE 0.020 WIDTH 0.080 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.020 SIDE 0.010 WIDTH 0.080 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.020 SIDE 0.020 WIDTH 0.120 ;
    ENCLOSURE CUTCLASS AYBAR BELOW END 0.030 SIDE 0.030 WIDTH 0.200 ;
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.002 SIDE 0.030 ;		 
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.030 SIDE 0.002 ;		 
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.007 SIDE 0.025 ;	     
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.025 SIDE 0.007 ;	     
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.020 SIDE 0.020 ;	     
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.005 SIDE 0.030 WIDTH 0.051 ;
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.030 SIDE 0.005 WIDTH 0.051 ;
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.010 SIDE 0.025 WIDTH 0.060 ;
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.025 SIDE 0.010 WIDTH 0.060 ;
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.020 SIDE 0.020 WIDTH 0.080 ;
    ENCLOSURE CUTCLASS AYBAR ABOVE END 0.030 SIDE 0.030 WIDTH 0.200 ; " ;	

# AY.EX.MLAST.2
    PROPERTY LEF58_EOLENCLOSURE "
    EOLENCLOSURE 0.105 CUTCLASS AY BELOW 0.020 MINLENGTH 0.021 ; " ; 
    
#AY.C.7 KEEPOUT rule. 
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C1 CUTCLASS AY NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C1 CUTCLASS AYBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;

# AY.S.CFIRST.1, AYBAR.S.CFIRST.1
  PROPERTY LEF58_SPACING "
	SPACING 0.015 LAYER C1 CUTCLASS AY CONCAVECORNER ;
	SPACING 0.02 LAYER C1 CUTCLASS AYBAR CONCAVECORNER ; " ;


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END AY



LAYER C1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.090 0.090 ;
  OFFSET 0 0 ;
  MINWIDTH 0.044 ;
  MAXWIDTH 4.100 ;                               # Cx.W.2
  WIDTH 0.044 ;
	      
# Cx.S.1       
    SPACING 0.046 ;

# Cx.SE.1
    MINSTEP 0.046 MAXEDGES 1 ; 

# Cx.A.1
    AREA 0.01100 ; 

# Cx.A.2
    PROPERTY LEF58_AREA "
        AREA 0.0243 EXCEPTEDGELENGTH 0.117 ; " ;
        
# Cx.A.3
    MINENCLOSEDAREA 0.16 ;
    
# Cx.S.2/3/5  (S.4 is overwritten by S.5 - slight pessimism)
    PROPERTY LEF58_SPACING "
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.046 ENDTOEND 0.072 MINLENGTH 0.021 TWOSIDES ;
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.023 PARALLELEDGE 0.115 WITHIN 0.050 TWOEDGES ; " ;
 
# Cx.S.6-11
    SPACINGTABLE
	PARALLELRUNLENGTH        0       0.197  0.422  0.566  1.349
        WIDTH   0                0.046   0.046  0.046  0.046  0.046
        WIDTH   0.081            0.046   0.054  0.054  0.054  0.054
        WIDTH   0.117            0.046   0.072  0.072  0.072  0.072
        WIDTH   0.144            0.046   0.090  0.090  0.090  0.090
        WIDTH   0.423            0.046   0.090  0.117  0.117  0.117
        WIDTH   0.567            0.046   0.090  0.117  0.135  0.135
        WIDTH   1.350            0.046   0.090  0.117  0.135  0.450 ;
           

#Ax.C.11-14 AY.C.12-15
 PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS AY 2  WIDTH 0.185 WITHIN 0.221 FROMBELOW ;
    MINIMUMCUT  CUTCLASS AYBAR 1 WIDTH 0.185 WITHIN 0.181 FROMBELOW ;
    MINIMUMCUT CUTCLASS AY 2 WIDTH 0.185 WITHIN 0.221 FROMBELOW LENGTH 0.185 WITHIN 1.401 ;
    MINIMUMCUT CUTCLASS AY 3  WIDTH 0.349 WITHIN 0.221 FROMBELOW ;
    MINIMUMCUT CUTCLASS AY 4  WIDTH 0.479 WITHIN 0.221 FROMBELOW ;
    MINIMUMCUT  CUTCLASS AYBAR 2  WIDTH 0.349 WITHIN 0.181 FROMBELOW ;
    MINIMUMCUT  CUTCLASS AYBAR 2  WIDTH 0.479 WITHIN 0.181 FROMBELOW ;
    MINIMUMCUT CUTCLASS Ax 2   WIDTH 0.193 WITHIN 0.217 FROMABOVE LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT  CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171 FROMABOVE LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT CUTCLASS Ax 2   WIDTH 0.193 WITHIN 0.217 FROMABOVE ;
    MINIMUMCUT CUTCLASS Ax 3   WIDTH 0.599 WITHIN 0.217 FROMABOVE ;
    MINIMUMCUT CUTCLASS Ax 4   WIDTH 0.899 WITHIN 0.217 FROMABOVE ;
    MINIMUMCUT  CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171 FROMABOVE ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.599 WITHIN 0.171 FROMABOVE ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.899 WITHIN 0.171 FROMABOVE ; " ; 



 PROPERTY LEF58_VOLTAGESPACING
   "VOLTAGESPACING
     1.32 0.046
     1.65 0.050
     1.98 0.060
     2.75 0.070
     3.63 0.100
     5.50 0.120
     7.70 0.150
     11.0 0.180
     16.5 0.200
     18.7 0.220 ; " ;


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END C1

LAYER A1
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS Ax    WIDTH 0.044000 CUTS 1 ;
    CUTCLASS AxBAR WIDTH 0.044000 LENGTH 0.090000 CUTS 2 ; " ; # Ax.LW.1, AxBAR.W.1 & AxBAR.L.1

  PROPERTY LEF58_SPACING "
    SPACING 0.134 CENTERTOCENTER ADJACENTCUTS 3 WITHIN 0.134 CUTCLASS Ax ; " ; # Ax.C.2

 PROPERTY LEF58_SPACINGTABLE "
 SPACINGTABLE
     CENTERTOCENTER Ax TO Ax
     CUTCLASS          Ax        AxBAR SIDE     AxBAR END      
     Ax          0.125  0.125  0.068  0.072  0.068  0.072 
     AxBAR SIDE  0.068  0.072  0.072  0.072  0.082  0.082 
     AxBAR END   0.068  0.072  0.082  0.082  0.092  0.092 ; " ; # Ax.S.1, Ax.S.AxBAR.S.1, AxBAR.S.1, Ax.S.AxBAR.S.2, AxBAR.S.2

#Ax.EX.Cx.1.or a/b/c
#Ax.EX.Cy.1.or a/b/c, Ax.EN.Cy.2
#AxBAR.EX.Cx.1.or a/b/c, Ax.EN.Cx.2,3
#AxBAR.EX.Cy.1.or a/b/c, Ax.EN.Cy.2,3
#
	PROPERTY LEF58_ENCLOSURE "
		ENCLOSURE CUTCLASS Ax 0.004000 0.020000 ;
		ENCLOSURE CUTCLASS Ax 0.018000 0.018000 ;
		ENCLOSURE CUTCLASS Ax BELOW 0.000000 0.025000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.000000 0.032000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.010000 0.020000 WIDTH 0.088000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.018000 0.018000 WIDTH 0.088000 ;

		ENCLOSURE CUTCLASS AxBAR END 0.036000 SIDE 0.000000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.018000 SIDE 0.018000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.009000 SIDE 0.027000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.027000 SIDE 0.009000 ;

		ENCLOSURE CUTCLASS AxBAR END 0.018000 SIDE 0.018000 WIDTH 0.084000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.023000 SIDE 0.023000 WIDTH 0.136000 ; " ;


    
#Ax.C.4 KEEPOUT rule. 
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C1 CUTCLASS Ax NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C2 CUTCLASS Ax NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C1 CUTCLASS AxBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C2 CUTCLASS AxBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;



  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END A1



LAYER C2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.090 0.090 ;
  OFFSET 0 0 ;
  MINWIDTH 0.044 ;
  MAXWIDTH 4.100 ;                               # Cx.W.2
  WIDTH 0.044 ;
	      
# Cx.S.1       
    SPACING 0.046 ;

# Cx.SE.1
    MINSTEP 0.046 MAXEDGES 1 ; 

# Cx.A.1
    AREA 0.01100 ; 

# Cx.A.2
    PROPERTY LEF58_AREA "
        AREA 0.0243 EXCEPTEDGELENGTH 0.117 ; " ;
        
# Cx.A.3
    MINENCLOSEDAREA 0.16 ;
    
# Cx.S.2/3/5  (S.4 is overwritten by S.5 - slight pessimism)
    PROPERTY LEF58_SPACING "
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.046 ENDTOEND 0.072 MINLENGTH 0.021 TWOSIDES ;
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.023 PARALLELEDGE 0.115 WITHIN 0.050 TWOEDGES ; " ;
 
# Cx.S.6-11
    SPACINGTABLE
	PARALLELRUNLENGTH        0       0.197  0.422  0.566  1.349
        WIDTH   0                0.046   0.046  0.046  0.046  0.046
        WIDTH   0.081            0.046   0.054  0.054  0.054  0.054
        WIDTH   0.117            0.046   0.072  0.072  0.072  0.072
        WIDTH   0.144            0.046   0.090  0.090  0.090  0.090
        WIDTH   0.423            0.046   0.090  0.117  0.117  0.117
        WIDTH   0.567            0.046   0.090  0.117  0.135  0.135
        WIDTH   1.350            0.046   0.090  0.117  0.135  0.450 ;
           

 PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS Ax 2    WIDTH 0.193 WITHIN 0.217  LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT   CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171  LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT CUTCLASS Ax 2   WIDTH 0.193 WITHIN 0.217  ;
    MINIMUMCUT CUTCLASS Ax 3   WIDTH 0.599 WITHIN 0.217  ;
    MINIMUMCUT CUTCLASS Ax 4   WIDTH 0.899 WITHIN 0.217  ; 
    MINIMUMCUT  CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171  ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.599 WITHIN 0.171  ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.899 WITHIN 0.171  ; " ;	     # Ax.C.11-14



 PROPERTY LEF58_VOLTAGESPACING
   "VOLTAGESPACING
     1.32 0.046
     1.65 0.050
     1.98 0.060
     2.75 0.070
     3.63 0.100
     5.50 0.120
     7.70 0.150
     11.0 0.180
     16.5 0.200
     18.7 0.220 ; " ;


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END C2

LAYER A2
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS Ax    WIDTH 0.044000 CUTS 1 ;
    CUTCLASS AxBAR WIDTH 0.044000 LENGTH 0.090000 CUTS 2 ; " ; # Ax.LW.1, AxBAR.W.1 & AxBAR.L.1

  PROPERTY LEF58_SPACING "
    SPACING 0.134 CENTERTOCENTER ADJACENTCUTS 3 WITHIN 0.134 CUTCLASS Ax ; " ; # Ax.C.2

 PROPERTY LEF58_SPACINGTABLE "
 SPACINGTABLE
     CENTERTOCENTER Ax TO Ax
     CUTCLASS          Ax        AxBAR SIDE     AxBAR END      
     Ax          0.125  0.125  0.068  0.072  0.068  0.072 
     AxBAR SIDE  0.068  0.072  0.072  0.072  0.082  0.082 
     AxBAR END   0.068  0.072  0.082  0.082  0.092  0.092 ; " ; # Ax.S.1, Ax.S.AxBAR.S.1, AxBAR.S.1, Ax.S.AxBAR.S.2, AxBAR.S.2

#Ax.EX.Cx.1.or a/b/c
#Ax.EX.Cy.1.or a/b/c, Ax.EN.Cy.2
#AxBAR.EX.Cx.1.or a/b/c, Ax.EN.Cx.2,3
#AxBAR.EX.Cy.1.or a/b/c, Ax.EN.Cy.2,3
#
	PROPERTY LEF58_ENCLOSURE "
		ENCLOSURE CUTCLASS Ax 0.004000 0.020000 ;
		ENCLOSURE CUTCLASS Ax 0.018000 0.018000 ;
		ENCLOSURE CUTCLASS Ax BELOW 0.000000 0.025000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.000000 0.032000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.010000 0.020000 WIDTH 0.088000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.018000 0.018000 WIDTH 0.088000 ;

		ENCLOSURE CUTCLASS AxBAR END 0.036000 SIDE 0.000000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.018000 SIDE 0.018000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.009000 SIDE 0.027000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.027000 SIDE 0.009000 ;

		ENCLOSURE CUTCLASS AxBAR END 0.018000 SIDE 0.018000 WIDTH 0.084000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.023000 SIDE 0.023000 WIDTH 0.136000 ; " ;


    
#Ax.C.4 KEEPOUT rule. 
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C2 CUTCLASS Ax NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C3 CUTCLASS Ax NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C2 CUTCLASS AxBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C3 CUTCLASS AxBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;



  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END A2



LAYER C3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.090 0.090 ;
  OFFSET 0 0 ;
  MINWIDTH 0.044 ;
  MAXWIDTH 4.100 ;                               # Cx.W.2
  WIDTH 0.044 ;
	      
# Cx.S.1       
    SPACING 0.046 ;

# Cx.SE.1
    MINSTEP 0.046 MAXEDGES 1 ; 

# Cx.A.1
    AREA 0.01100 ; 

# Cx.A.2
    PROPERTY LEF58_AREA "
        AREA 0.0243 EXCEPTEDGELENGTH 0.117 ; " ;
        
# Cx.A.3
    MINENCLOSEDAREA 0.16 ;
    
# Cx.S.2/3/5  (S.4 is overwritten by S.5 - slight pessimism)
    PROPERTY LEF58_SPACING "
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.046 ENDTOEND 0.072 MINLENGTH 0.021 TWOSIDES ;
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.023 PARALLELEDGE 0.115 WITHIN 0.050 TWOEDGES ; " ;
 
# Cx.S.6-11
    SPACINGTABLE
	PARALLELRUNLENGTH        0       0.197  0.422  0.566  1.349
        WIDTH   0                0.046   0.046  0.046  0.046  0.046
        WIDTH   0.081            0.046   0.054  0.054  0.054  0.054
        WIDTH   0.117            0.046   0.072  0.072  0.072  0.072
        WIDTH   0.144            0.046   0.090  0.090  0.090  0.090
        WIDTH   0.423            0.046   0.090  0.117  0.117  0.117
        WIDTH   0.567            0.046   0.090  0.117  0.135  0.135
        WIDTH   1.350            0.046   0.090  0.117  0.135  0.450 ;
           

 PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS Ax 2    WIDTH 0.193 WITHIN 0.217  LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT   CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171  LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT CUTCLASS Ax 2   WIDTH 0.193 WITHIN 0.217  ;
    MINIMUMCUT CUTCLASS Ax 3   WIDTH 0.599 WITHIN 0.217  ;
    MINIMUMCUT CUTCLASS Ax 4   WIDTH 0.899 WITHIN 0.217  ; 
    MINIMUMCUT  CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171  ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.599 WITHIN 0.171  ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.899 WITHIN 0.171  ; " ;	     # Ax.C.11-14



 PROPERTY LEF58_VOLTAGESPACING
   "VOLTAGESPACING
     1.32 0.046
     1.65 0.050
     1.98 0.060
     2.75 0.070
     3.63 0.100
     5.50 0.120
     7.70 0.150
     11.0 0.180
     16.5 0.200
     18.7 0.220 ; " ;


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END C3

LAYER A3
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS Ax    WIDTH 0.044000 CUTS 1 ;
    CUTCLASS AxBAR WIDTH 0.044000 LENGTH 0.090000 CUTS 2 ; " ; # Ax.LW.1, AxBAR.W.1 & AxBAR.L.1

  PROPERTY LEF58_SPACING "
    SPACING 0.134 CENTERTOCENTER ADJACENTCUTS 3 WITHIN 0.134 CUTCLASS Ax ; " ; # Ax.C.2

 PROPERTY LEF58_SPACINGTABLE "
 SPACINGTABLE
     CENTERTOCENTER Ax TO Ax
     CUTCLASS          Ax        AxBAR SIDE     AxBAR END      
     Ax          0.125  0.125  0.068  0.072  0.068  0.072 
     AxBAR SIDE  0.068  0.072  0.072  0.072  0.082  0.082 
     AxBAR END   0.068  0.072  0.082  0.082  0.092  0.092 ; " ; # Ax.S.1, Ax.S.AxBAR.S.1, AxBAR.S.1, Ax.S.AxBAR.S.2, AxBAR.S.2

#Ax.EX.Cx.1.or a/b/c
#Ax.EX.Cy.1.or a/b/c, Ax.EN.Cy.2
#AxBAR.EX.Cx.1.or a/b/c, Ax.EN.Cx.2,3
#AxBAR.EX.Cy.1.or a/b/c, Ax.EN.Cy.2,3
#
	PROPERTY LEF58_ENCLOSURE "
		ENCLOSURE CUTCLASS Ax 0.004000 0.020000 ;
		ENCLOSURE CUTCLASS Ax 0.018000 0.018000 ;
		ENCLOSURE CUTCLASS Ax BELOW 0.000000 0.025000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.000000 0.032000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.010000 0.020000 WIDTH 0.088000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.018000 0.018000 WIDTH 0.088000 ;

		ENCLOSURE CUTCLASS AxBAR END 0.036000 SIDE 0.000000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.018000 SIDE 0.018000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.009000 SIDE 0.027000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.027000 SIDE 0.009000 ;

		ENCLOSURE CUTCLASS AxBAR END 0.018000 SIDE 0.018000 WIDTH 0.084000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.023000 SIDE 0.023000 WIDTH 0.136000 ; " ;


    
#Ax.C.4 KEEPOUT rule. 
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C3 CUTCLASS Ax NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C4 CUTCLASS Ax NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C3 CUTCLASS AxBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C4 CUTCLASS AxBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;



  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END A3



LAYER C4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.090 0.090 ;
  OFFSET 0 0 ;
  MINWIDTH 0.044 ;
  MAXWIDTH 4.100 ;                               # Cx.W.2
  WIDTH 0.044 ;
	      
# Cx.S.1       
    SPACING 0.046 ;

# Cx.SE.1
    MINSTEP 0.046 MAXEDGES 1 ; 

# Cx.A.1
    AREA 0.01100 ; 

# Cx.A.2
    PROPERTY LEF58_AREA "
        AREA 0.0243 EXCEPTEDGELENGTH 0.117 ; " ;
        
# Cx.A.3
    MINENCLOSEDAREA 0.16 ;
    
# Cx.S.2/3/5  (S.4 is overwritten by S.5 - slight pessimism)
    PROPERTY LEF58_SPACING "
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.046 ENDTOEND 0.072 MINLENGTH 0.021 TWOSIDES ;
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.023 PARALLELEDGE 0.115 WITHIN 0.050 TWOEDGES ; " ;
 
# Cx.S.6-11
    SPACINGTABLE
	PARALLELRUNLENGTH        0       0.197  0.422  0.566  1.349
        WIDTH   0                0.046   0.046  0.046  0.046  0.046
        WIDTH   0.081            0.046   0.054  0.054  0.054  0.054
        WIDTH   0.117            0.046   0.072  0.072  0.072  0.072
        WIDTH   0.144            0.046   0.090  0.090  0.090  0.090
        WIDTH   0.423            0.046   0.090  0.117  0.117  0.117
        WIDTH   0.567            0.046   0.090  0.117  0.135  0.135
        WIDTH   1.350            0.046   0.090  0.117  0.135  0.450 ;
           

 PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS Ax 2    WIDTH 0.193 WITHIN 0.217  LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT   CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171  LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT CUTCLASS Ax 2   WIDTH 0.193 WITHIN 0.217  ;
    MINIMUMCUT CUTCLASS Ax 3   WIDTH 0.599 WITHIN 0.217  ;
    MINIMUMCUT CUTCLASS Ax 4   WIDTH 0.899 WITHIN 0.217  ; 
    MINIMUMCUT  CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171  ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.599 WITHIN 0.171  ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.899 WITHIN 0.171  ; " ;	     # Ax.C.11-14



 PROPERTY LEF58_VOLTAGESPACING
   "VOLTAGESPACING
     1.32 0.046
     1.65 0.050
     1.98 0.060
     2.75 0.070
     3.63 0.100
     5.50 0.120
     7.70 0.150
     11.0 0.180
     16.5 0.200
     18.7 0.220 ; " ;


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END C4

LAYER A4
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS Ax    WIDTH 0.044000 CUTS 1 ;
    CUTCLASS AxBAR WIDTH 0.044000 LENGTH 0.090000 CUTS 2 ; " ; # Ax.LW.1, AxBAR.W.1 & AxBAR.L.1

  PROPERTY LEF58_SPACING "
    SPACING 0.134 CENTERTOCENTER ADJACENTCUTS 3 WITHIN 0.134 CUTCLASS Ax ; " ; # Ax.C.2

 PROPERTY LEF58_SPACINGTABLE "
 SPACINGTABLE
     CENTERTOCENTER Ax TO Ax
     CUTCLASS          Ax        AxBAR SIDE     AxBAR END      
     Ax          0.125  0.125  0.068  0.072  0.068  0.072 
     AxBAR SIDE  0.068  0.072  0.072  0.072  0.082  0.082 
     AxBAR END   0.068  0.072  0.082  0.082  0.092  0.092 ; " ; # Ax.S.1, Ax.S.AxBAR.S.1, AxBAR.S.1, Ax.S.AxBAR.S.2, AxBAR.S.2

#Ax.EX.Cx.1.or a/b/c
#Ax.EX.Cy.1.or a/b/c, Ax.EN.Cy.2
#AxBAR.EX.Cx.1.or a/b/c, Ax.EN.Cx.2,3
#AxBAR.EX.Cy.1.or a/b/c, Ax.EN.Cy.2,3
#
	PROPERTY LEF58_ENCLOSURE "
		ENCLOSURE CUTCLASS Ax 0.004000 0.020000 ;
		ENCLOSURE CUTCLASS Ax 0.018000 0.018000 ;
		ENCLOSURE CUTCLASS Ax BELOW 0.000000 0.025000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.000000 0.032000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.010000 0.020000 WIDTH 0.088000 ;
		ENCLOSURE CUTCLASS Ax ABOVE 0.018000 0.018000 WIDTH 0.088000 ;

		ENCLOSURE CUTCLASS AxBAR END 0.036000 SIDE 0.000000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.018000 SIDE 0.018000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.009000 SIDE 0.027000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.027000 SIDE 0.009000 ;

		ENCLOSURE CUTCLASS AxBAR END 0.018000 SIDE 0.018000 WIDTH 0.084000 ;
		ENCLOSURE CUTCLASS AxBAR END 0.023000 SIDE 0.023000 WIDTH 0.136000 ; " ;


    
#Ax.C.4 KEEPOUT rule. 
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C4 CUTCLASS Ax NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C5 CUTCLASS Ax NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C4 CUTCLASS AxBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;
 PROPERTY LEF58_SPACING "SPACING 0.035 LAYER C5 CUTCLASS AxBAR NONEOLCONVEXCORNER 0.061 MINLENGTH 0.021 ;" ;



  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END A4



LAYER C5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.090 0.090 ;
  OFFSET 0 0 ;
  MINWIDTH 0.044 ;
  MAXWIDTH 4.100 ;                               # Cx.W.2
  WIDTH 0.044 ;
	      
# Cx.S.1       
    SPACING 0.046 ;

# Cx.SE.1
    MINSTEP 0.046 MAXEDGES 1 ; 

# Cx.A.1
    AREA 0.01100 ; 

# Cx.A.2
    PROPERTY LEF58_AREA "
        AREA 0.0243 EXCEPTEDGELENGTH 0.117 ; " ;
        
# Cx.A.3
    MINENCLOSEDAREA 0.16 ;
    
# Cx.S.2/3/5  (S.4 is overwritten by S.5 - slight pessimism)
    PROPERTY LEF58_SPACING "
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.046 ENDTOEND 0.072 MINLENGTH 0.021 TWOSIDES ;
      SPACING 0.063 ENDOFLINE 0.101 WITHIN 0.023 PARALLELEDGE 0.115 WITHIN 0.050 TWOEDGES ; " ;
 
# Cx.S.6-11
    SPACINGTABLE
	PARALLELRUNLENGTH        0       0.197  0.422  0.566  1.349
        WIDTH   0                0.046   0.046  0.046  0.046  0.046
        WIDTH   0.081            0.046   0.054  0.054  0.054  0.054
        WIDTH   0.117            0.046   0.072  0.072  0.072  0.072
        WIDTH   0.144            0.046   0.090  0.090  0.090  0.090
        WIDTH   0.423            0.046   0.090  0.117  0.117  0.117
        WIDTH   0.567            0.046   0.090  0.117  0.135  0.135
        WIDTH   1.350            0.046   0.090  0.117  0.135  0.450 ;
           

 PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS Ax 2    WIDTH 0.193 WITHIN 0.217 FROMBELOW LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT   CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171 FROMBELOW LENGTH 0.193 WITHIN 1.401 ;
    MINIMUMCUT CUTCLASS Ax 2   WIDTH 0.193 WITHIN 0.217 FROMBELOW ;
    MINIMUMCUT CUTCLASS Ax 3   WIDTH 0.599 WITHIN 0.217 FROMBELOW ;
    MINIMUMCUT CUTCLASS Ax 4   WIDTH 0.899 WITHIN 0.217 FROMBELOW ; 
    MINIMUMCUT  CUTCLASS AxBAR 1  WIDTH 0.193 WITHIN 0.171 FROMBELOW ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.599 WITHIN 0.171 FROMBELOW ;
    MINIMUMCUT  CUTCLASS AxBAR 2  WIDTH 0.899 WITHIN 0.171 FROMBELOW ; " ;    # Ax.C.11-14, no YS.C. rules defined



 PROPERTY LEF58_VOLTAGESPACING
   "VOLTAGESPACING
     1.32 0.046
     1.65 0.050
     1.98 0.060
     2.75 0.070
     3.63 0.100
     5.50 0.120
     7.70 0.150
     11.0 0.180
     16.5 0.200
     18.7 0.220 ; " ;


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END C5

LAYER YS
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS YS       WIDTH 0.414 ; " ;            # YS.LW.1
  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
    CUTCLASS    YS 
    YS          0.486 0.486 ; " ;                  # table values: noPRL, PRL, YS.S.2
  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
    SAMENET
    CUTCLASS    YS 
    YS          0.396 0.396 ; " ;                  # table values: noPRL, PRL, YS.S.1 
  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS YS 0.018 0.072 ; " ;        # YS.EN/EX....
  
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END YS

LAYER JA
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH  0.90 ; 
  OFFSET 0.0 0.0 ;                          # user input, floorplan/stdcell dependent  
  WIDTH 0.450 ;                             # Jx.W.1
  MINWIDTH 0.450 ;                          # Jx.W.1

  SPACINGTABLE TWOWIDTHS         					# Jx.S.2 - 8
		###	width=	0.000	1.500	4.500	
		###	prl=	none	1.500	4.500
		###	-------------------------------------
    WIDTH 0.000 	        0.450	0.585   1.350
    WIDTH 1.500 PRL 1.500       0.585   0.585   1.350
    WIDTH 4.500 PRL 4.500	1.350	1.350	1.350 ;

  AREA 0.810 ;                              # Jx.A.1
  MAXWIDTH 10.8   ;                         # Jx.W.2
  MINENCLOSEDAREA 0.810 ;                   # Jx.A.2


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END JA


LAYER JV
  TYPE CUT ;

    PROPERTY LEF58_CUTCLASS "
                CUTCLASS JV    WIDTH 1.20 CUTS 1 ; " ;	# JV.LW.1

    PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
        CUTCLASS          JV     
        JV             1.20  1.20  ; " ;	  # JV.S.1, JVBAR.S.1, JVBAR.S.JV.1


    PROPERTY LEF58_ENCLOSURE "
        ENCLOSURE CUTCLASS JV BELOW 0.30 0.60 ;
        ENCLOSURE CUTCLASS JV ABOVE 0.60 0.30 ; " ;  # JV.EX.JLAST.2, JV.EN.QA.2
 

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END JV

# 30x layer - only basic rules are supported
LAYER QA
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 2.4 2.4 ;
  OFFSET 0.0 0.0 ;
  WIDTH 1.2 ;                              # Qx.W.1  
  MINWIDTH 1.2 ;                           # Qx.W.1
  SPACINGTABLE TWOWIDTHS         	   # Qx.S.1/2/3  PRL only for S.3 valid!
		###	width=	0.000	6.000    6.000 
		###	prl=	none	none     6.000
		###	-------------------------------
    WIDTH 0.000 	        1.200	1.800    1.800
    WIDTH 6.000 	        1.800   1.800    1.800 
    WIDTH 6.000  PRL 6.000      1.800   1.800    2.400 ;
  AREA 2 ;                                 # Qx.A.1
  MINENCLOSEDAREA 2 ;	                   # Qx.A.2
  MAXWIDTH 18 ;                            # Qx.W.2

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END QA


LAYER JW
  TYPE CUT ;

    PROPERTY LEF58_CUTCLASS "
                CUTCLASS JW    WIDTH 1.20 CUTS 1 ; " ;	# JW.LW.1

    PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
        CUTCLASS          JW     
        JW             1.20  1.20  ; " ;	  # JW.S.1


    PROPERTY LEF58_ENCLOSURE "
        ENCLOSURE CUTCLASS JW BELOW 0.30 0.60 ;
        ENCLOSURE CUTCLASS JW ABOVE 0.60 0.30 ; " ;  # JW.EN.QA.2, JW.EX.Qx.1
 

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 20.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 5.0 ;
  ANTENNAGATEPLUSDIFF 5.0 ;

END JW

# 30x layer - only basic rules are supported
LAYER QB
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 2.4 2.4 ;
  OFFSET 0.0 0.0 ;
  WIDTH 1.2 ;                              # Qx.W.1  
  MINWIDTH 1.2 ;                           # Qx.W.1
  SPACINGTABLE TWOWIDTHS         	   # Qx.S.1/2/3  PRL only for S.3 valid!
		###	width=	0.000	6.000    6.000 
		###	prl=	none	none     6.000
		###	-------------------------------
    WIDTH 0.000 	        1.200	1.800    1.800
    WIDTH 6.000 	        1.800   1.800    1.800 
    WIDTH 6.000  PRL 6.000      1.800   1.800    2.400 ;
  AREA 2 ;                                 # Qx.A.1
  MINENCLOSEDAREA 2 ;	                   # Qx.A.2
  MAXWIDTH 18 ;                            # Qx.W.2

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END QB


LAYER VV
  TYPE CUT ;

    PROPERTY LEF58_CUTCLASS "
                CUTCLASS VV    WIDTH 2.70 CUTS 1 ; " ;	# VV.LW.1

# VV.S.1
    PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
        CUTCLASS          VV
        VV             1.80  1.80 ; " ;	# VV.S.1

# VV.EN.LM.1 VV.EN.LB.1 
    PROPERTY LEF58_ENCLOSURE "

        ENCLOSURE CUTCLASS VV BELOW 0.450 0.450 ;
        ENCLOSURE CUTCLASS VV ABOVE 0.450 0.450 ; " ;	# VV.EN.LM.1, VV.EN.LB.1



  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAAREAFACTOR 10000 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 20000 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAAREAFACTOR 10000 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 20000 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAAREAFACTOR 10000 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 20000 ;" ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAAREAFACTOR 10000 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 20000 ;" ;

END VV

LAYER LB
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 3.6 3.6 ;
  WIDTH 1.8 ;
  SPACING 1.8 ;
  MAXWIDTH 100 ;      # dummy

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;
  ANTENNAMODEL OXIDE4 ;
  ANTENNADIFFAREARATIO 500.0 ;
  ANTENNAGATEPLUSDIFF 2.0 ;

END LB



LAYER OVERLAP
TYPE OVERLAP ;
END OVERLAP


#################################################

#################################################


#------------------------------------------------------------
#  V1 VIA SECTION 
#------------------------------------------------------------
 VIA VIA01_0_30_0_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_0_30_0_30_HH_V1
 
 VIA VIA01_0_30_0_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_0_30_0_30_HV_V1
 
 VIA VIA01 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01
 
 VIA VIA01_I DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_I
 
 VIA VIA01_0_30_3_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_0_30_3_30_HH_V1
 
 VIA VIA01_0_30_3_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_0_30_3_30_HV_V1
 
 VIA VIA01_0_30_3_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_0_30_3_30_VH_V1
 
 VIA VIA01_0_30_3_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_0_30_3_30_VV_V1
 
 VIA VIA01_0_30_5_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_0_30_5_30_HH_V1
 
 VIA VIA01_0_30_5_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_0_30_5_30_HV_V1
 
 VIA VIA01_0_30_5_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_0_30_5_30_VH_V1
 
 VIA VIA01_0_30_5_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_0_30_5_30_VV_V1
 
 VIA VIA01_0_30_7_25_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_0_30_7_25_HH_V1
 
 VIA VIA01_0_30_7_25_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_0_30_7_25_HV_V1
 
 VIA VIA01_0_30_7_25_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_0_30_7_25_VH_V1
 
 VIA VIA01_0_30_7_25_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_0_30_7_25_VV_V1
 
 VIA VIA01_0_30_10_25_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_0_30_10_25_HH_V1
 
 VIA VIA01_0_30_10_25_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_0_30_10_25_HV_V1
 
 VIA VIA01_0_30_10_25_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_0_30_10_25_VH_V1
 
 VIA VIA01_0_30_10_25_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_0_30_10_25_VV_V1
 
 VIA VIA01_0_30_20_20_HX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_0_30_20_20_HX_V1
 
 VIA VIA01_0_30_20_20_VX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_0_30_20_20_VX_V1
 
 VIA VIA01_0_30_25_25_HX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_0_30_25_25_HX_V1
 
 VIA VIA01_0_30_25_25_VX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_0_30_25_25_VX_V1
 
 VIA VIA01_5_30_0_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_5_30_0_30_HH_V1
 
 VIA VIA01_5_30_0_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_5_30_0_30_HV_V1
 
 VIA VIA01_5_30_0_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_5_30_0_30_VH_V1
 
 VIA VIA01_5_30_0_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_5_30_0_30_VV_V1
 
 VIA VIA01_5_30_3_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_5_30_3_30_HH_V1
 
 VIA VIA01_5_30_3_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_5_30_3_30_HV_V1
 
 VIA VIA01_5_30_3_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_5_30_3_30_VH_V1
 
 VIA VIA01_5_30_3_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_5_30_3_30_VV_V1
 
 VIA VIA01_5_30_5_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_5_30_5_30_HH_V1
 
 VIA VIA01_5_30_5_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_5_30_5_30_HV_V1
 
 VIA VIA01_5_30_5_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_5_30_5_30_VH_V1
 
 VIA VIA01_5_30_5_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_5_30_5_30_VV_V1
 
 VIA VIA01_5_30_7_25_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_5_30_7_25_HH_V1
 
 VIA VIA01_5_30_7_25_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_5_30_7_25_HV_V1
 
 VIA VIA01_5_30_7_25_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_5_30_7_25_VH_V1
 
 VIA VIA01_5_30_7_25_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_5_30_7_25_VV_V1
 
 VIA VIA01_5_30_10_25_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_5_30_10_25_HH_V1
 
 VIA VIA01_5_30_10_25_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_5_30_10_25_HV_V1
 
 VIA VIA01_5_30_10_25_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_5_30_10_25_VH_V1
 
 VIA VIA01_5_30_10_25_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_5_30_10_25_VV_V1
 
 VIA VIA01_5_30_20_20_HX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_5_30_20_20_HX_V1
 
 VIA VIA01_5_30_20_20_VX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_5_30_20_20_VX_V1
 
 VIA VIA01_5_30_25_25_HX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_5_30_25_25_HX_V1
 
 VIA VIA01_5_30_25_25_VX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_5_30_25_25_VX_V1
 
 VIA VIA01_10_20_0_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_10_20_0_30_HH_V1
 
 VIA VIA01_10_20_0_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_10_20_0_30_HV_V1
 
 VIA VIA01_10_20_0_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_10_20_0_30_VH_V1
 
 VIA VIA01_10_20_0_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_10_20_0_30_VV_V1
 
 VIA VIA01_10_20_3_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_10_20_3_30_HH_V1
 
 VIA VIA01_10_20_3_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_10_20_3_30_HV_V1
 
 VIA VIA01_10_20_3_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_10_20_3_30_VH_V1
 
 VIA VIA01_10_20_3_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_10_20_3_30_VV_V1
 
 VIA VIA01_10_20_5_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_10_20_5_30_HH_V1
 
 VIA VIA01_10_20_5_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_10_20_5_30_HV_V1
 
 VIA VIA01_10_20_5_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_10_20_5_30_VH_V1
 
 VIA VIA01_10_20_5_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_10_20_5_30_VV_V1
 
 VIA VIA01_10_20_7_25_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_10_20_7_25_HH_V1
 
 VIA VIA01_10_20_7_25_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_10_20_7_25_HV_V1
 
 VIA VIA01_10_20_7_25_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_10_20_7_25_VH_V1
 
 VIA VIA01_10_20_7_25_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_10_20_7_25_VV_V1
 
 VIA VIA01_10_20_10_25_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_10_20_10_25_HH_V1
 
 VIA VIA01_10_20_10_25_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_10_20_10_25_HV_V1
 
 VIA VIA01_10_20_10_25_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_10_20_10_25_VH_V1
 
 VIA VIA01_10_20_10_25_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_10_20_10_25_VV_V1
 
 VIA VIA01_10_20_20_20_HX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_10_20_20_20_HX_V1
 
 VIA VIA01_10_20_20_20_VX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_10_20_20_20_VX_V1
 
 VIA VIA01_10_20_25_25_HX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.030 0.040 0.030 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_10_20_25_25_HX_V1
 
 VIA VIA01_10_20_25_25_VX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_10_20_25_25_VX_V1
 
 VIA VIA01_7_25_0_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_7_25_0_30_HH_V1
 
 VIA VIA01_7_25_0_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_7_25_0_30_HV_V1
 
 VIA VIA01_7_25_0_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_7_25_0_30_VH_V1
 
 VIA VIA01_7_25_0_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_7_25_0_30_VV_V1
 
 VIA VIA01_7_25_3_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_7_25_3_30_HH_V1
 
 VIA VIA01_7_25_3_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_7_25_3_30_HV_V1
 
 VIA VIA01_7_25_3_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_7_25_3_30_VH_V1
 
 VIA VIA01_7_25_3_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_7_25_3_30_VV_V1
 
 VIA VIA01_7_25_5_30_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_7_25_5_30_HH_V1
 
 VIA VIA01_7_25_5_30_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_7_25_5_30_HV_V1
 
 VIA VIA01_7_25_5_30_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_7_25_5_30_VH_V1
 
 VIA VIA01_7_25_5_30_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_7_25_5_30_VV_V1
 
 VIA VIA01_7_25_7_25_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_7_25_7_25_HH_V1
 
 VIA VIA01_7_25_7_25_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_7_25_7_25_HV_V1
 
 VIA VIA01_7_25_7_25_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_7_25_7_25_VH_V1
 
 VIA VIA01_7_25_7_25_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_7_25_7_25_VV_V1
 
 VIA VIA01_7_25_10_25_HH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_7_25_10_25_HH_V1
 
 VIA VIA01_7_25_10_25_HV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_7_25_10_25_HV_V1
 
 VIA VIA01_7_25_10_25_VH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_7_25_10_25_VH_V1
 
 VIA VIA01_7_25_10_25_VV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_7_25_10_25_VV_V1
 
 VIA VIA01_7_25_20_20_HX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_7_25_20_20_HX_V1
 
 VIA VIA01_7_25_20_20_VX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_7_25_20_20_VX_V1
 
 VIA VIA01_7_25_25_25_HX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_7_25_25_25_HX_V1
 
 VIA VIA01_7_25_25_25_VX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_7_25_25_25_VX_V1
 
 VIA VIA01_20_20_0_30_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_20_20_0_30_XH_V1
 
 VIA VIA01_20_20_0_30_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_20_20_0_30_XV_V1
 
 VIA VIA01_20_20_3_30_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_20_20_3_30_XH_V1
 
 VIA VIA01_20_20_3_30_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_20_20_3_30_XV_V1
 
 VIA VIA01_20_20_5_30_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_20_20_5_30_XH_V1
 
 VIA VIA01_20_20_5_30_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_20_20_5_30_XV_V1
 
 VIA VIA01_20_20_7_25_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_20_20_7_25_XH_V1
 
 VIA VIA01_20_20_7_25_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_20_20_7_25_XV_V1
 
 VIA VIA01_20_20_10_25_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_20_20_10_25_XH_V1
 
 VIA VIA01_20_20_10_25_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_20_20_10_25_XV_V1
 
 VIA VIA01_20_20_20_20_XX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_20_20_20_20_XX_V1
 
 VIA VIA01_20_20_25_25_XX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_20_20_25_25_XX_V1
 
 VIA VIA01_25_25_0_30_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 END VIA01_25_25_0_30_XH_V1
 
 VIA VIA01_25_25_0_30_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 END VIA01_25_25_0_30_XV_V1
 
 VIA VIA01_25_25_3_30_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 END VIA01_25_25_3_30_XH_V1
 
 VIA VIA01_25_25_3_30_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.023 -0.050 0.023 0.050 ;
 END VIA01_25_25_3_30_XV_V1
 
 VIA VIA01_25_25_5_30_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 END VIA01_25_25_5_30_XH_V1
 
 VIA VIA01_25_25_5_30_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 END VIA01_25_25_5_30_XV_V1
 
 VIA VIA01_25_25_7_25_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 END VIA01_25_25_7_25_XH_V1
 
 VIA VIA01_25_25_7_25_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 END VIA01_25_25_7_25_XV_V1
 
 VIA VIA01_25_25_10_25_XH_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 END VIA01_25_25_10_25_XH_V1
 
 VIA VIA01_25_25_10_25_XV_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.030 -0.045 0.030 0.045 ;
 END VIA01_25_25_10_25_XV_V1
 
 VIA VIA01_25_25_20_20_XX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA01_25_25_20_20_XX_V1
 
 VIA VIA01_25_25_25_25_XX_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 LAYER M2 ;
 RECT -0.045 -0.045 0.045 0.045 ;
 END VIA01_25_25_25_25_XX_V1
 
 VIA VIA01_BAR_V_0_30_0_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_BAR_V_0_30_0_30_V1
 
 VIA VIA01_BAR_V_0_30_3_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 LAYER M2 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 END VIA01_BAR_V_0_30_3_30_V1
 
 VIA VIA01_BAR_V_0_30_5_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 LAYER M2 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 END VIA01_BAR_V_0_30_5_30_V1
 
 VIA VIA01_BAR_V_0_30_7_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 LAYER M2 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 END VIA01_BAR_V_0_30_7_25_V1
 
 VIA VIA01_BAR_V_0_30_10_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 LAYER M2 ;
 RECT -0.030 -0.065 0.030 0.065 ;
 END VIA01_BAR_V_0_30_10_25_V1
 
 VIA VIA01_BAR_V_0_30_20_20_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 LAYER M2 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 END VIA01_BAR_V_0_30_20_20_V1
 
 VIA VIA01_BAR_V_0_30_30_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 LAYER M2 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 END VIA01_BAR_V_0_30_30_30_V1
 
 VIA VIA01_BAR_V_3_30_0_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_BAR_V_3_30_0_30_V1
 
 VIA VIA01_BAR_V_3_30_3_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 LAYER M2 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 END VIA01_BAR_V_3_30_3_30_V1
 
 VIA VIA01_BAR_V_3_30_5_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 LAYER M2 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 END VIA01_BAR_V_3_30_5_30_V1
 
 VIA VIA01_BAR_V_3_30_7_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 LAYER M2 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 END VIA01_BAR_V_3_30_7_25_V1
 
 VIA VIA01_BAR_V_3_30_10_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 LAYER M2 ;
 RECT -0.030 -0.065 0.030 0.065 ;
 END VIA01_BAR_V_3_30_10_25_V1
 
 VIA VIA01_BAR_V_3_30_20_20_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 LAYER M2 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 END VIA01_BAR_V_3_30_20_20_V1
 
 VIA VIA01_BAR_V_3_30_30_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 LAYER M2 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 END VIA01_BAR_V_3_30_30_30_V1
 
 VIA VIA01_BAR_V_5_30_0_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_BAR_V_5_30_0_30_V1
 
 VIA VIA01_BAR_V_5_30_3_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 LAYER M2 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 END VIA01_BAR_V_5_30_3_30_V1
 
 VIA VIA01_BAR_V_5_30_5_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 LAYER M2 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 END VIA01_BAR_V_5_30_5_30_V1
 
 VIA VIA01_BAR_V_5_30_7_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 LAYER M2 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 END VIA01_BAR_V_5_30_7_25_V1
 
 VIA VIA01_BAR_V_5_30_10_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 LAYER M2 ;
 RECT -0.030 -0.065 0.030 0.065 ;
 END VIA01_BAR_V_5_30_10_25_V1
 
 VIA VIA01_BAR_V_5_30_20_20_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 LAYER M2 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 END VIA01_BAR_V_5_30_20_20_V1
 
 VIA VIA01_BAR_V_5_30_30_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 LAYER M2 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 END VIA01_BAR_V_5_30_30_30_V1
 
 VIA VIA01_BAR_V_7_25_0_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_BAR_V_7_25_0_30_V1
 
 VIA VIA01_BAR_V_7_25_3_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 LAYER M2 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 END VIA01_BAR_V_7_25_3_30_V1
 
 VIA VIA01_BAR_V_7_25_5_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 LAYER M2 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 END VIA01_BAR_V_7_25_5_30_V1
 
 VIA VIA01_BAR_V_7_25_7_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 LAYER M2 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 END VIA01_BAR_V_7_25_7_25_V1
 
 VIA VIA01_BAR_V_7_25_10_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 LAYER M2 ;
 RECT -0.030 -0.065 0.030 0.065 ;
 END VIA01_BAR_V_7_25_10_25_V1
 
 VIA VIA01_BAR_V_7_25_20_20_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 LAYER M2 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 END VIA01_BAR_V_7_25_20_20_V1
 
 VIA VIA01_BAR_V_7_25_30_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 LAYER M2 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 END VIA01_BAR_V_7_25_30_30_V1
 
 VIA VIA01_BAR_V_10_20_0_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.030 -0.060 0.030 0.060 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_BAR_V_10_20_0_30_V1
 
 VIA VIA01_BAR_V_10_20_3_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.030 -0.060 0.030 0.060 ;
 LAYER M2 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 END VIA01_BAR_V_10_20_3_30_V1
 
 VIA VIA01_BAR_V_10_20_5_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.030 -0.060 0.030 0.060 ;
 LAYER M2 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 END VIA01_BAR_V_10_20_5_30_V1
 
 VIA VIA01_BAR_V_10_20_7_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.030 -0.060 0.030 0.060 ;
 LAYER M2 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 END VIA01_BAR_V_10_20_7_25_V1
 
 VIA VIA01_BAR_V_10_20_10_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.030 -0.060 0.030 0.060 ;
 LAYER M2 ;
 RECT -0.030 -0.065 0.030 0.065 ;
 END VIA01_BAR_V_10_20_10_25_V1
 
 VIA VIA01_BAR_V_10_20_20_20_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.030 -0.060 0.030 0.060 ;
 LAYER M2 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 END VIA01_BAR_V_10_20_20_20_V1
 
 VIA VIA01_BAR_V_10_20_30_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.030 -0.060 0.030 0.060 ;
 LAYER M2 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 END VIA01_BAR_V_10_20_30_30_V1
 
 VIA VIA01_BAR_V_20_20_0_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_BAR_V_20_20_0_30_V1
 
 VIA VIA01_BAR_V_20_20_3_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 LAYER M2 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 END VIA01_BAR_V_20_20_3_30_V1
 
 VIA VIA01_BAR_V_20_20_5_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 LAYER M2 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 END VIA01_BAR_V_20_20_5_30_V1
 
 VIA VIA01_BAR_V_20_20_7_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 LAYER M2 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 END VIA01_BAR_V_20_20_7_25_V1
 
 VIA VIA01_BAR_V_20_20_10_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 LAYER M2 ;
 RECT -0.030 -0.065 0.030 0.065 ;
 END VIA01_BAR_V_20_20_10_25_V1
 
 VIA VIA01_BAR_V_20_20_20_20_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 LAYER M2 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 END VIA01_BAR_V_20_20_20_20_V1
 
 VIA VIA01_BAR_V_20_20_30_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 LAYER M2 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 END VIA01_BAR_V_20_20_30_30_V1
 
 VIA VIA01_BAR_V_30_30_0_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_BAR_V_30_30_0_30_V1
 
 VIA VIA01_BAR_V_30_30_3_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 LAYER M2 ;
 RECT -0.023 -0.070 0.023 0.070 ;
 END VIA01_BAR_V_30_30_3_30_V1
 
 VIA VIA01_BAR_V_30_30_5_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 LAYER M2 ;
 RECT -0.025 -0.070 0.025 0.070 ;
 END VIA01_BAR_V_30_30_5_30_V1
 
 VIA VIA01_BAR_V_30_30_7_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 LAYER M2 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 END VIA01_BAR_V_30_30_7_25_V1
 
 VIA VIA01_BAR_V_30_30_10_25_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 LAYER M2 ;
 RECT -0.030 -0.065 0.030 0.065 ;
 END VIA01_BAR_V_30_30_10_25_V1
 
 VIA VIA01_BAR_V_30_30_20_20_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 LAYER M2 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 END VIA01_BAR_V_30_30_20_20_V1
 
 VIA VIA01_BAR_V_30_30_30_30_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M1 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 LAYER M2 ;
 RECT -0.050 -0.070 0.050 0.070 ;
 END VIA01_BAR_V_30_30_30_30_V1
 
 VIA VIA01_BAR_H_0_30_0_30_V1_LW DEFAULT
 LAYER V1 ;
 RECT -0.090 -0.020 -0.010 0.020 ;
 LAYER M1 ;
 RECT -0.120 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.120 -0.020 0.020 0.020 ;
 END VIA01_BAR_H_0_30_0_30_V1_LW
 
 VIA VIA01_BAR_H_0_30_0_30_V1_LE DEFAULT
 LAYER V1 ;
 RECT 0.010 -0.020 0.090 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.020 0.120 0.020 ;
 LAYER M2 ;
 RECT -0.020 -0.020 0.120 0.020 ;
 END VIA01_BAR_H_0_30_0_30_V1_LE
 
 VIA VIA01_BAR_H_10_20_0_30_V1_LW DEFAULT
 LAYER V1 ;
 RECT -0.080 -0.020 0.000 0.020 ;
 LAYER M1 ;
 RECT -0.100 -0.030 0.020 0.030 ;
 LAYER M2 ;
 RECT -0.110 -0.020 0.030 0.020 ;
 END VIA01_BAR_H_10_20_0_30_V1_LW
 
 VIA VIA01_BAR_H_10_20_0_30_V1_LE DEFAULT
 LAYER V1 ;
 RECT 0.000 -0.020 0.080 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.030 0.100 0.030 ;
 LAYER M2 ;
 RECT -0.030 -0.020 0.110 0.020 ;
 END VIA01_BAR_H_10_20_0_30_V1_LE
 
 VIA VIA01_BAR_V_10_20_0_30_V1_LW DEFAULT
 LAYER V1 ;
 RECT -0.030 -0.040 0.010 0.040 ;
 LAYER M1 ;
 RECT -0.040 -0.060 0.020 0.060 ;
 LAYER M2 ;
 RECT -0.030 -0.070 0.010 0.070 ;
 END VIA01_BAR_V_10_20_0_30_V1_LW
 
 VIA VIA01_BAR_V_10_20_0_30_V1_LE DEFAULT
 LAYER V1 ;
 RECT -0.010 -0.040 0.030 0.040 ;
 LAYER M1 ;
 RECT -0.020 -0.060 0.040 0.060 ;
 LAYER M2 ;
 RECT -0.010 -0.070 0.030 0.070 ;
 END VIA01_BAR_V_10_20_0_30_V1_LE
 
 VIA VIA01_BAR_V_0_30_0_30_V1_UN DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.090 0.020 -0.010 ;
 LAYER M1 ;
 RECT -0.020 -0.120 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.020 -0.120 0.020 0.020 ;
 END VIA01_BAR_V_0_30_0_30_V1_UN
 
 VIA VIA01_BAR_V_0_30_0_30_V1_US DEFAULT
 LAYER V1 ;
 RECT -0.020 0.010 0.020 0.090 ;
 LAYER M1 ;
 RECT -0.020 -0.020 0.020 0.120 ;
 LAYER M2 ;
 RECT -0.020 -0.020 0.020 0.120 ;
 END VIA01_BAR_V_0_30_0_30_V1_US
 
 VIA VIA01_BAR_V_10_20_0_30_V1_UN DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.090 0.020 -0.010 ;
 LAYER M1 ;
 RECT -0.030 -0.110 0.030 0.010 ;
 LAYER M2 ;
 RECT -0.020 -0.120 0.020 0.020 ;
 END VIA01_BAR_V_10_20_0_30_V1_UN
 
 VIA VIA01_BAR_V_10_20_0_30_V1_US DEFAULT
 LAYER V1 ;
 RECT -0.020 0.010 0.020 0.090 ;
 LAYER M1 ;
 RECT -0.030 -0.010 0.030 0.110 ;
 LAYER M2 ;
 RECT -0.020 -0.020 0.020 0.120 ;
 END VIA01_BAR_V_10_20_0_30_V1_US
 
 VIA VIA01_0_30_0_35_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.055 -0.020 0.055 0.020 ;
 END VIA01_0_30_0_35_VH_V1_R
 
 VIA VIA01_0_30_0_35_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.055 0.020 0.055 ;
 END VIA01_0_30_0_35_VV_V1_R
 
 VIA VIA01_0_30_0_40_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.060 -0.020 0.060 0.020 ;
 END VIA01_0_30_0_40_VH_V1_R
 
 VIA VIA01_0_30_0_40_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.060 0.020 0.060 ;
 END VIA01_0_30_0_40_VV_V1_R
 
 VIA VIA01_0_30_0_50_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 END VIA01_0_30_0_50_VH_V1_R
 
 VIA VIA01_0_30_0_50_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_0_30_0_50_VV_V1_R
 
 VIA VIA01_0_30_0_60_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.080 -0.020 0.080 0.020 ;
 END VIA01_0_30_0_60_VH_V1_R
 
 VIA VIA01_0_30_0_60_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.020 -0.050 0.020 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.080 0.020 0.080 ;
 END VIA01_0_30_0_60_VV_V1_R
 
 VIA VIA01_5_30_0_35_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.055 -0.020 0.055 0.020 ;
 END VIA01_5_30_0_35_VH_V1_R
 
 VIA VIA01_5_30_0_35_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.055 0.020 0.055 ;
 END VIA01_5_30_0_35_VV_V1_R
 
 VIA VIA01_5_30_0_40_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.060 -0.020 0.060 0.020 ;
 END VIA01_5_30_0_40_VH_V1_R
 
 VIA VIA01_5_30_0_40_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.060 0.020 0.060 ;
 END VIA01_5_30_0_40_VV_V1_R
 
 VIA VIA01_5_30_0_50_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 END VIA01_5_30_0_50_VH_V1_R
 
 VIA VIA01_5_30_0_50_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_5_30_0_50_VV_V1_R
 
 VIA VIA01_5_30_0_60_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.080 -0.020 0.080 0.020 ;
 END VIA01_5_30_0_60_VH_V1_R
 
 VIA VIA01_5_30_0_60_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.025 -0.050 0.025 0.050 ;
 LAYER M2 ;
 RECT -0.020 -0.080 0.020 0.080 ;
 END VIA01_5_30_0_60_VV_V1_R
 
 VIA VIA01_10_20_0_35_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.055 -0.020 0.055 0.020 ;
 END VIA01_10_20_0_35_VH_V1_R
 
 VIA VIA01_10_20_0_35_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.020 -0.055 0.020 0.055 ;
 END VIA01_10_20_0_35_VV_V1_R
 
 VIA VIA01_10_20_0_40_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.060 -0.020 0.060 0.020 ;
 END VIA01_10_20_0_40_VH_V1_R
 
 VIA VIA01_10_20_0_40_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.020 -0.060 0.020 0.060 ;
 END VIA01_10_20_0_40_VV_V1_R
 
 VIA VIA01_10_20_0_50_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 END VIA01_10_20_0_50_VH_V1_R
 
 VIA VIA01_10_20_0_50_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_10_20_0_50_VV_V1_R
 
 VIA VIA01_10_20_0_60_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.080 -0.020 0.080 0.020 ;
 END VIA01_10_20_0_60_VH_V1_R
 
 VIA VIA01_10_20_0_60_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.030 -0.040 0.030 0.040 ;
 LAYER M2 ;
 RECT -0.020 -0.080 0.020 0.080 ;
 END VIA01_10_20_0_60_VV_V1_R
 
 VIA VIA01_7_25_0_35_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.055 -0.020 0.055 0.020 ;
 END VIA01_7_25_0_35_VH_V1_R
 
 VIA VIA01_7_25_0_35_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.020 -0.055 0.020 0.055 ;
 END VIA01_7_25_0_35_VV_V1_R
 
 VIA VIA01_7_25_0_40_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.060 -0.020 0.060 0.020 ;
 END VIA01_7_25_0_40_VH_V1_R
 
 VIA VIA01_7_25_0_40_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.020 -0.060 0.020 0.060 ;
 END VIA01_7_25_0_40_VV_V1_R
 
 VIA VIA01_7_25_0_50_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 END VIA01_7_25_0_50_VH_V1_R
 
 VIA VIA01_7_25_0_50_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.020 -0.070 0.020 0.070 ;
 END VIA01_7_25_0_50_VV_V1_R
 
 VIA VIA01_7_25_0_60_VH_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.080 -0.020 0.080 0.020 ;
 END VIA01_7_25_0_60_VH_V1_R
 
 VIA VIA01_7_25_0_60_VV_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M1 ;
 RECT -0.027 -0.045 0.027 0.045 ;
 LAYER M2 ;
 RECT -0.020 -0.080 0.020 0.080 ;
 END VIA01_7_25_0_60_VV_V1_R
 
 VIA VIA01_BAR_H_7_25_0_37_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M1 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 LAYER M2 ;
 RECT -0.077 -0.020 0.077 0.020 ;
 END VIA01_BAR_H_7_25_0_37_V1_R
 
 VIA VIA01_BAR_H_10_20_0_37_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M1 ;
 RECT -0.060 -0.030 0.060 0.030 ;
 LAYER M2 ;
 RECT -0.077 -0.020 0.077 0.020 ;
 END VIA01_BAR_H_10_20_0_37_V1_R
 
 VIA VIA01_BAR_H_20_20_0_37_V1_R DEFAULT
 LAYER V1 ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M1 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 LAYER M2 ;
 RECT -0.077 -0.020 0.077 0.020 ;
 END VIA01_BAR_H_20_20_0_37_V1_R
 
 VIA VIA01_20_20_20_20_VH_2CUT_H_V1 DEFAULT
 LAYER V1 ;
 RECT -0.078 -0.020 -0.038 0.020 ;
 RECT 0.038 -0.020 0.078 0.020 ;
 LAYER M1 ;
 RECT -0.098 -0.040 0.098 0.040 ;
 LAYER M2 ;
 RECT -0.098 -0.040 0.098 0.040 ;
 END VIA01_20_20_20_20_VH_2CUT_H_V1
 
 VIA VIA01_20_20_20_20_VH_2CUT_V_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.078 0.020 -0.038 ;
 RECT -0.020 0.038 0.020 0.078 ;
 LAYER M1 ;
 RECT -0.040 -0.098 0.040 0.098 ;
 LAYER M2 ;
 RECT -0.040 -0.098 0.040 0.098 ;
 END VIA01_20_20_20_20_VH_2CUT_V_V1
 
 VIA VIA01_0_30_20_20_VH_2CUT_V_V1 DEFAULT
 LAYER V1 ;
 RECT -0.020 -0.078 0.020 -0.038 ;
 RECT -0.020 0.038 0.020 0.078 ;
 LAYER M1 ;
 RECT -0.020 -0.108 0.020 0.108 ;
 LAYER M2 ;
 RECT -0.040 -0.098 0.040 0.098 ;
 END VIA01_0_30_20_20_VH_2CUT_V_V1
 
 VIA VIA01_20_20_20_20_XX_4CUT_V1 DEFAULT
 LAYER V1 ;
 RECT -0.085 -0.085 -0.045 -0.045 ;
 RECT 0.045 -0.085 0.085 -0.045 ;
 RECT -0.085 0.045 -0.045 0.085 ;
 RECT 0.045 0.045 0.085 0.085 ;
 LAYER M1 ;
 RECT -0.105 -0.105 0.105 0.105 ;
 LAYER M2 ;
 RECT -0.105 -0.105 0.105 0.105 ;
 END VIA01_20_20_20_20_XX_4CUT_V1
 
VIARULE VIA01_GEN_0_30_0_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.000 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.000 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_0_30_0_30_VH_V1 

VIARULE VIA01_GEN_0_30_3_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.000 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.003 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_0_30_3_30_VH_V1 

VIARULE VIA01_GEN_0_30_5_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.000 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_0_30_5_30_VH_V1 

VIARULE VIA01_GEN_0_30_10_25_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.000 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_0_30_10_25_VH_V1 

VIARULE VIA01_GEN_0_30_20_20_VX_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.000 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_0_30_20_20_VX_V1 

VIARULE VIA01_GEN_0_30_30_30_VX_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.000 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.030 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_0_30_30_30_VX_V1 

VIARULE VIA01_GEN_5_30_0_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.000 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_5_30_0_30_VH_V1 

VIARULE VIA01_GEN_5_30_3_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.003 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_5_30_3_30_VH_V1 

VIARULE VIA01_GEN_5_30_5_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_5_30_5_30_VH_V1 

VIARULE VIA01_GEN_5_30_10_25_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_5_30_10_25_VH_V1 

VIARULE VIA01_GEN_5_30_20_20_VX_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_5_30_20_20_VX_V1 

VIARULE VIA01_GEN_5_30_30_30_VX_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.030 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_5_30_30_30_VX_V1 

VIARULE VIA01_GEN_10_20_0_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.010 0.020 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.000 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_10_20_0_30_VH_V1 

VIARULE VIA01_GEN_10_20_3_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.010 0.020 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.003 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_10_20_3_30_VH_V1 

VIARULE VIA01_GEN_10_20_5_30_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.010 0.020 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_10_20_5_30_VH_V1 

VIARULE VIA01_GEN_10_20_10_25_VH_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.010 0.020 ;
  LAYER M2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_10_20_10_25_VH_V1 

VIARULE VIA01_GEN_10_20_20_20_VX_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.010 0.020 ;
  LAYER M2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_10_20_20_20_VX_V1 

VIARULE VIA01_GEN_10_20_30_30_VX_V1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.010 0.020 ;
  LAYER M2 ;
    ENCLOSURE 0.030 0.030 ;
  LAYER V1 ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.115 ;
END  VIA01_GEN_10_20_30_30_VX_V1 

#------------------------------------------------------------
#  AY VIA SECTION 
#------------------------------------------------------------
 VIA VIA02_0_30_2_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA02_0_30_2_34_HH_AY
 
 VIA VIA02 DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA02
 
 VIA VIA02_0_30_5_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.054 -0.025 0.054 0.025 ;
 END VIA02_0_30_5_34_HH_AY
 
 VIA VIA02_0_30_5_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.025 -0.054 0.025 0.054 ;
 END VIA02_0_30_5_34_HV_AY
 
 VIA VIA02_0_30_7_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.050 -0.027 0.050 0.027 ;
 END VIA02_0_30_7_30_HH_AY
 
 VIA VIA02_0_30_7_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.027 -0.050 0.027 0.050 ;
 END VIA02_0_30_7_30_HV_AY
 
 VIA VIA02_0_30_10_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.050 -0.030 0.050 0.030 ;
 END VIA02_0_30_10_30_HH_AY
 
 VIA VIA02_0_30_10_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.030 -0.050 0.030 0.050 ;
 END VIA02_0_30_10_30_HV_AY
 
 VIA VIA02_0_30_20_20_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA02_0_30_20_20_HX_AY
 
 VIA VIA02_0_30_30_30_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 END VIA02_0_30_30_30_HX_AY
 
 VIA VIA02_3_30_2_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA02_3_30_2_34_HH_AY
 
 VIA VIA02_3_30_2_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA02_3_30_2_34_HV_AY
 
 VIA VIA02_3_30_5_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.054 -0.025 0.054 0.025 ;
 END VIA02_3_30_5_34_HH_AY
 
 VIA VIA02_3_30_5_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.025 -0.054 0.025 0.054 ;
 END VIA02_3_30_5_34_HV_AY
 
 VIA VIA02_3_30_7_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.050 -0.027 0.050 0.027 ;
 END VIA02_3_30_7_30_HH_AY
 
 VIA VIA02_3_30_7_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.027 -0.050 0.027 0.050 ;
 END VIA02_3_30_7_30_HV_AY
 
 VIA VIA02_3_30_10_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.050 -0.030 0.050 0.030 ;
 END VIA02_3_30_10_30_HH_AY
 
 VIA VIA02_3_30_10_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.030 -0.050 0.030 0.050 ;
 END VIA02_3_30_10_30_HV_AY
 
 VIA VIA02_3_30_20_20_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA02_3_30_20_20_HX_AY
 
 VIA VIA02_3_30_30_30_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 END VIA02_3_30_30_30_HX_AY
 
 VIA VIA02_5_30_2_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA02_5_30_2_34_HH_AY
 
 VIA VIA02_5_30_2_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA02_5_30_2_34_HV_AY
 
 VIA VIA02_5_30_5_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.054 -0.025 0.054 0.025 ;
 END VIA02_5_30_5_34_HH_AY
 
 VIA VIA02_5_30_5_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.025 -0.054 0.025 0.054 ;
 END VIA02_5_30_5_34_HV_AY
 
 VIA VIA02_5_30_7_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.050 -0.027 0.050 0.027 ;
 END VIA02_5_30_7_30_HH_AY
 
 VIA VIA02_5_30_7_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.027 -0.050 0.027 0.050 ;
 END VIA02_5_30_7_30_HV_AY
 
 VIA VIA02_5_30_10_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.050 -0.030 0.050 0.030 ;
 END VIA02_5_30_10_30_HH_AY
 
 VIA VIA02_5_30_10_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.030 -0.050 0.030 0.050 ;
 END VIA02_5_30_10_30_HV_AY
 
 VIA VIA02_5_30_20_20_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA02_5_30_20_20_HX_AY
 
 VIA VIA02_5_30_30_30_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 END VIA02_5_30_30_30_HX_AY
 
 VIA VIA02_7_25_2_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA02_7_25_2_34_HH_AY
 
 VIA VIA02_7_25_2_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA02_7_25_2_34_HV_AY
 
 VIA VIA02_7_25_5_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.054 -0.025 0.054 0.025 ;
 END VIA02_7_25_5_34_HH_AY
 
 VIA VIA02_7_25_5_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.025 -0.054 0.025 0.054 ;
 END VIA02_7_25_5_34_HV_AY
 
 VIA VIA02_7_25_7_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.050 -0.027 0.050 0.027 ;
 END VIA02_7_25_7_30_HH_AY
 
 VIA VIA02_7_25_7_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.027 -0.050 0.027 0.050 ;
 END VIA02_7_25_7_30_HV_AY
 
 VIA VIA02_7_25_10_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.050 -0.030 0.050 0.030 ;
 END VIA02_7_25_10_30_HH_AY
 
 VIA VIA02_7_25_10_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.030 -0.050 0.030 0.050 ;
 END VIA02_7_25_10_30_HV_AY
 
 VIA VIA02_7_25_20_20_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA02_7_25_20_20_HX_AY
 
 VIA VIA02_7_25_30_30_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 END VIA02_7_25_30_30_HX_AY
 
 VIA VIA02_10_25_2_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA02_10_25_2_34_HH_AY
 
 VIA VIA02_10_25_2_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA02_10_25_2_34_HV_AY
 
 VIA VIA02_10_25_5_34_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.054 -0.025 0.054 0.025 ;
 END VIA02_10_25_5_34_HH_AY
 
 VIA VIA02_10_25_5_34_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.025 -0.054 0.025 0.054 ;
 END VIA02_10_25_5_34_HV_AY
 
 VIA VIA02_10_25_7_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.050 -0.027 0.050 0.027 ;
 END VIA02_10_25_7_30_HH_AY
 
 VIA VIA02_10_25_7_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.027 -0.050 0.027 0.050 ;
 END VIA02_10_25_7_30_HV_AY
 
 VIA VIA02_10_25_10_30_HH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.050 -0.030 0.050 0.030 ;
 END VIA02_10_25_10_30_HH_AY
 
 VIA VIA02_10_25_10_30_HV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.030 -0.050 0.030 0.050 ;
 END VIA02_10_25_10_30_HV_AY
 
 VIA VIA02_10_25_20_20_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA02_10_25_20_20_HX_AY
 
 VIA VIA02_10_25_30_30_HX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 END VIA02_10_25_30_30_HX_AY
 
 VIA VIA02_20_20_2_34_XH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA02_20_20_2_34_XH_AY
 
 VIA VIA02_20_20_2_34_XV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA02_20_20_2_34_XV_AY
 
 VIA VIA02_20_20_5_34_XH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.054 -0.025 0.054 0.025 ;
 END VIA02_20_20_5_34_XH_AY
 
 VIA VIA02_20_20_5_34_XV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.025 -0.054 0.025 0.054 ;
 END VIA02_20_20_5_34_XV_AY
 
 VIA VIA02_20_20_7_30_XH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.050 -0.027 0.050 0.027 ;
 END VIA02_20_20_7_30_XH_AY
 
 VIA VIA02_20_20_7_30_XV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.027 -0.050 0.027 0.050 ;
 END VIA02_20_20_7_30_XV_AY
 
 VIA VIA02_20_20_10_30_XH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.050 -0.030 0.050 0.030 ;
 END VIA02_20_20_10_30_XH_AY
 
 VIA VIA02_20_20_10_30_XV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.030 -0.050 0.030 0.050 ;
 END VIA02_20_20_10_30_XV_AY
 
 VIA VIA02_20_20_20_20_XX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA02_20_20_20_20_XX_AY
 
 VIA VIA02_20_20_30_30_XX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 END VIA02_20_20_30_30_XX_AY
 
 VIA VIA02_30_30_2_34_XH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA02_30_30_2_34_XH_AY
 
 VIA VIA02_30_30_2_34_XV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA02_30_30_2_34_XV_AY
 
 VIA VIA02_30_30_5_34_XH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.054 -0.025 0.054 0.025 ;
 END VIA02_30_30_5_34_XH_AY
 
 VIA VIA02_30_30_5_34_XV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.025 -0.054 0.025 0.054 ;
 END VIA02_30_30_5_34_XV_AY
 
 VIA VIA02_30_30_7_30_XH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.050 -0.027 0.050 0.027 ;
 END VIA02_30_30_7_30_XH_AY
 
 VIA VIA02_30_30_7_30_XV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.027 -0.050 0.027 0.050 ;
 END VIA02_30_30_7_30_XV_AY
 
 VIA VIA02_30_30_10_30_XH_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.050 -0.030 0.050 0.030 ;
 END VIA02_30_30_10_30_XH_AY
 
 VIA VIA02_30_30_10_30_XV_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.030 -0.050 0.030 0.050 ;
 END VIA02_30_30_10_30_XV_AY
 
 VIA VIA02_30_30_20_20_XX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA02_30_30_20_20_XX_AY
 
 VIA VIA02_30_30_30_30_XX_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 END VIA02_30_30_30_30_XX_AY
 
 VIA VIA02_BAR_H_0_30_2_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 LAYER C1 ;
 RECT -0.070 -0.022 0.070 0.022 ;
 END VIA02_BAR_H_0_30_2_30_AY
 
 VIA VIA02_BAR_H_0_30_5_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 LAYER C1 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 END VIA02_BAR_H_0_30_5_30_AY
 
 VIA VIA02_BAR_H_0_30_7_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 LAYER C1 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 END VIA02_BAR_H_0_30_7_25_AY
 
 VIA VIA02_BAR_H_0_30_10_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 LAYER C1 ;
 RECT -0.065 -0.030 0.065 0.030 ;
 END VIA02_BAR_H_0_30_10_25_AY
 
 VIA VIA02_BAR_H_0_30_20_20_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 LAYER C1 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 END VIA02_BAR_H_0_30_20_20_AY
 
 VIA VIA02_BAR_H_0_30_30_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 LAYER C1 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 END VIA02_BAR_H_0_30_30_30_AY
 
 VIA VIA02_BAR_H_3_30_2_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.023 0.070 0.023 ;
 LAYER C1 ;
 RECT -0.070 -0.022 0.070 0.022 ;
 END VIA02_BAR_H_3_30_2_30_AY
 
 VIA VIA02_BAR_H_3_30_5_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.023 0.070 0.023 ;
 LAYER C1 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 END VIA02_BAR_H_3_30_5_30_AY
 
 VIA VIA02_BAR_H_3_30_7_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.023 0.070 0.023 ;
 LAYER C1 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 END VIA02_BAR_H_3_30_7_25_AY
 
 VIA VIA02_BAR_H_3_30_10_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.023 0.070 0.023 ;
 LAYER C1 ;
 RECT -0.065 -0.030 0.065 0.030 ;
 END VIA02_BAR_H_3_30_10_25_AY
 
 VIA VIA02_BAR_H_3_30_20_20_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.023 0.070 0.023 ;
 LAYER C1 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 END VIA02_BAR_H_3_30_20_20_AY
 
 VIA VIA02_BAR_H_3_30_30_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.023 0.070 0.023 ;
 LAYER C1 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 END VIA02_BAR_H_3_30_30_30_AY
 
 VIA VIA02_BAR_H_7_25_2_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 LAYER C1 ;
 RECT -0.070 -0.022 0.070 0.022 ;
 END VIA02_BAR_H_7_25_2_30_AY
 
 VIA VIA02_BAR_H_7_25_5_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 LAYER C1 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 END VIA02_BAR_H_7_25_5_30_AY
 
 VIA VIA02_BAR_H_7_25_7_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 LAYER C1 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 END VIA02_BAR_H_7_25_7_25_AY
 
 VIA VIA02_BAR_H_7_25_10_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 LAYER C1 ;
 RECT -0.065 -0.030 0.065 0.030 ;
 END VIA02_BAR_H_7_25_10_25_AY
 
 VIA VIA02_BAR_H_7_25_20_20_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 LAYER C1 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 END VIA02_BAR_H_7_25_20_20_AY
 
 VIA VIA02_BAR_H_7_25_30_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 LAYER C1 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 END VIA02_BAR_H_7_25_30_30_AY
 
 VIA VIA02_BAR_H_5_30_2_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 LAYER C1 ;
 RECT -0.070 -0.022 0.070 0.022 ;
 END VIA02_BAR_H_5_30_2_30_AY
 
 VIA VIA02_BAR_H_5_30_5_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 LAYER C1 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 END VIA02_BAR_H_5_30_5_30_AY
 
 VIA VIA02_BAR_H_5_30_7_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 LAYER C1 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 END VIA02_BAR_H_5_30_7_25_AY
 
 VIA VIA02_BAR_H_5_30_10_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 LAYER C1 ;
 RECT -0.065 -0.030 0.065 0.030 ;
 END VIA02_BAR_H_5_30_10_25_AY
 
 VIA VIA02_BAR_H_5_30_20_20_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 LAYER C1 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 END VIA02_BAR_H_5_30_20_20_AY
 
 VIA VIA02_BAR_H_5_30_30_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 LAYER C1 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 END VIA02_BAR_H_5_30_30_30_AY
 
 VIA VIA02_BAR_H_10_20_2_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.030 0.060 0.030 ;
 LAYER C1 ;
 RECT -0.070 -0.022 0.070 0.022 ;
 END VIA02_BAR_H_10_20_2_30_AY
 
 VIA VIA02_BAR_H_10_20_5_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.030 0.060 0.030 ;
 LAYER C1 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 END VIA02_BAR_H_10_20_5_30_AY
 
 VIA VIA02_BAR_H_10_20_7_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.030 0.060 0.030 ;
 LAYER C1 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 END VIA02_BAR_H_10_20_7_25_AY
 
 VIA VIA02_BAR_H_10_20_10_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.030 0.060 0.030 ;
 LAYER C1 ;
 RECT -0.065 -0.030 0.065 0.030 ;
 END VIA02_BAR_H_10_20_10_25_AY
 
 VIA VIA02_BAR_H_10_20_20_20_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.030 0.060 0.030 ;
 LAYER C1 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 END VIA02_BAR_H_10_20_20_20_AY
 
 VIA VIA02_BAR_H_10_20_30_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.030 0.060 0.030 ;
 LAYER C1 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 END VIA02_BAR_H_10_20_30_30_AY
 
 VIA VIA02_BAR_H_20_20_2_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 LAYER C1 ;
 RECT -0.070 -0.022 0.070 0.022 ;
 END VIA02_BAR_H_20_20_2_30_AY
 
 VIA VIA02_BAR_H_20_20_5_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 LAYER C1 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 END VIA02_BAR_H_20_20_5_30_AY
 
 VIA VIA02_BAR_H_20_20_7_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 LAYER C1 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 END VIA02_BAR_H_20_20_7_25_AY
 
 VIA VIA02_BAR_H_20_20_10_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 LAYER C1 ;
 RECT -0.065 -0.030 0.065 0.030 ;
 END VIA02_BAR_H_20_20_10_25_AY
 
 VIA VIA02_BAR_H_20_20_20_20_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 LAYER C1 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 END VIA02_BAR_H_20_20_20_20_AY
 
 VIA VIA02_BAR_H_20_20_30_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 LAYER C1 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 END VIA02_BAR_H_20_20_30_30_AY
 
 VIA VIA02_BAR_H_30_30_2_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 LAYER C1 ;
 RECT -0.070 -0.022 0.070 0.022 ;
 END VIA02_BAR_H_30_30_2_30_AY
 
 VIA VIA02_BAR_H_30_30_5_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 LAYER C1 ;
 RECT -0.070 -0.025 0.070 0.025 ;
 END VIA02_BAR_H_30_30_5_30_AY
 
 VIA VIA02_BAR_H_30_30_7_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 LAYER C1 ;
 RECT -0.065 -0.027 0.065 0.027 ;
 END VIA02_BAR_H_30_30_7_25_AY
 
 VIA VIA02_BAR_H_30_30_10_25_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 LAYER C1 ;
 RECT -0.065 -0.030 0.065 0.030 ;
 END VIA02_BAR_H_30_30_10_25_AY
 
 VIA VIA02_BAR_H_30_30_20_20_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 LAYER C1 ;
 RECT -0.060 -0.040 0.060 0.040 ;
 END VIA02_BAR_H_30_30_20_20_AY
 
 VIA VIA02_BAR_H_30_30_30_30_AY DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 LAYER C1 ;
 RECT -0.070 -0.050 0.070 0.050 ;
 END VIA02_BAR_H_30_30_30_30_AY
 
 VIA VIA02_BAR_V_20_10_2_30_AY_LN DEFAULT
 LAYER AY ;
 RECT -0.020 -0.070 0.020 0.010 ;
 LAYER M2 ;
 RECT -0.040 -0.080 0.040 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.100 0.022 0.040 ;
 END VIA02_BAR_V_20_10_2_30_AY_LN
 
 VIA VIA02_BAR_V_20_10_2_30_AY_LS DEFAULT
 LAYER AY ;
 RECT -0.020 -0.010 0.020 0.070 ;
 LAYER M2 ;
 RECT -0.040 -0.020 0.040 0.080 ;
 LAYER C1 ;
 RECT -0.022 -0.040 0.022 0.100 ;
 END VIA02_BAR_V_20_10_2_30_AY_LS
 
 VIA VIA02_0_30_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_0_30_2_53_HH_AY_R
 
 VIA VIA02_0_30_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_0_30_2_53_HV_AY_R
 
 VIA VIA02_0_30_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_0_30_2_63_HH_AY_R
 
 VIA VIA02_0_30_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.020 0.050 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_0_30_2_63_HV_AY_R
 
 VIA VIA02_3_30_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_3_30_2_53_HH_AY_R
 
 VIA VIA02_3_30_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_3_30_2_53_HV_AY_R
 
 VIA VIA02_3_30_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_3_30_2_63_HH_AY_R
 
 VIA VIA02_3_30_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.023 0.050 0.023 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_3_30_2_63_HV_AY_R
 
 VIA VIA02_5_30_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_5_30_2_53_HH_AY_R
 
 VIA VIA02_5_30_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_5_30_2_53_HV_AY_R
 
 VIA VIA02_5_30_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_5_30_2_63_HH_AY_R
 
 VIA VIA02_5_30_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.025 0.050 0.025 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_5_30_2_63_HV_AY_R
 
 VIA VIA02_7_25_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_7_25_2_53_HH_AY_R
 
 VIA VIA02_7_25_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_7_25_2_53_HV_AY_R
 
 VIA VIA02_7_25_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_7_25_2_63_HH_AY_R
 
 VIA VIA02_7_25_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.027 0.045 0.027 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_7_25_2_63_HV_AY_R
 
 VIA VIA02_10_25_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_10_25_2_53_HH_AY_R
 
 VIA VIA02_10_25_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_10_25_2_53_HV_AY_R
 
 VIA VIA02_10_25_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_10_25_2_63_HH_AY_R
 
 VIA VIA02_10_25_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.045 -0.030 0.045 0.030 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_10_25_2_63_HV_AY_R
 
 VIA VIA02_20_20_2_53_XH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_20_20_2_53_XH_AY_R
 
 VIA VIA02_20_20_2_53_XV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_20_20_2_53_XV_AY_R
 
 VIA VIA02_20_20_2_63_XH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_20_20_2_63_XH_AY_R
 
 VIA VIA02_20_20_2_63_XV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_20_20_2_63_XV_AY_R
 
 VIA VIA02_30_30_2_53_XH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_30_30_2_53_XH_AY_R
 
 VIA VIA02_30_30_2_53_XV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_30_30_2_53_XV_AY_R
 
 VIA VIA02_30_30_2_63_XH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_30_30_2_63_XH_AY_R
 
 VIA VIA02_30_30_2_63_XV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.050 -0.050 0.050 0.050 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_30_30_2_63_XV_AY_R
 
 VIA VIA02_0_35_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.055 -0.020 0.055 0.020 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_0_35_2_53_HH_AY_R
 
 VIA VIA02_0_35_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.055 -0.020 0.055 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_0_35_2_53_HV_AY_R
 
 VIA VIA02_0_35_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.055 -0.020 0.055 0.020 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_0_35_2_63_HH_AY_R
 
 VIA VIA02_0_35_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.055 -0.020 0.055 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_0_35_2_63_HV_AY_R
 
 VIA VIA02_0_40_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.020 0.060 0.020 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_0_40_2_53_HH_AY_R
 
 VIA VIA02_0_40_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.020 0.060 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_0_40_2_53_HV_AY_R
 
 VIA VIA02_0_40_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.020 0.060 0.020 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_0_40_2_63_HH_AY_R
 
 VIA VIA02_0_40_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.060 -0.020 0.060 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_0_40_2_63_HV_AY_R
 
 VIA VIA02_0_53_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.073 -0.020 0.073 0.020 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_0_53_2_53_HH_AY_R
 
 VIA VIA02_0_53_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.073 -0.020 0.073 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_0_53_2_53_HV_AY_R
 
 VIA VIA02_0_53_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.073 -0.020 0.073 0.020 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_0_53_2_63_HH_AY_R
 
 VIA VIA02_0_53_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.073 -0.020 0.073 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_0_53_2_63_HV_AY_R
 
 VIA VIA02_0_63_2_53_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.083 -0.020 0.083 0.020 ;
 LAYER C1 ;
 RECT -0.073 -0.022 0.073 0.022 ;
 END VIA02_0_63_2_53_HH_AY_R
 
 VIA VIA02_0_63_2_53_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.083 -0.020 0.083 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.073 0.022 0.073 ;
 END VIA02_0_63_2_53_HV_AY_R
 
 VIA VIA02_0_63_2_63_HH_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.083 -0.020 0.083 0.020 ;
 LAYER C1 ;
 RECT -0.083 -0.022 0.083 0.022 ;
 END VIA02_0_63_2_63_HH_AY_R
 
 VIA VIA02_0_63_2_63_HV_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.020 0.020 0.020 ;
 LAYER M2 ;
 RECT -0.083 -0.020 0.083 0.020 ;
 LAYER C1 ;
 RECT -0.022 -0.083 0.022 0.083 ;
 END VIA02_0_63_2_63_HV_AY_R
 
 VIA VIA02_BAR_V_7_25_2_55_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M2 ;
 RECT -0.027 -0.065 0.027 0.065 ;
 LAYER C1 ;
 RECT -0.022 -0.095 0.022 0.095 ;
 END VIA02_BAR_V_7_25_2_55_AY_R
 
 VIA VIA02_BAR_V_10_25_2_55_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M2 ;
 RECT -0.030 -0.065 0.030 0.065 ;
 LAYER C1 ;
 RECT -0.022 -0.095 0.022 0.095 ;
 END VIA02_BAR_V_10_25_2_55_AY_R
 
 VIA VIA02_BAR_V_20_20_2_55_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.040 0.020 0.040 ;
 LAYER M2 ;
 RECT -0.040 -0.060 0.040 0.060 ;
 LAYER C1 ;
 RECT -0.022 -0.095 0.022 0.095 ;
 END VIA02_BAR_V_20_20_2_55_AY_R
 
 VIA VIA02_BAR_H_0_30_22_22_AY_R DEFAULT
 LAYER AY ;
 RECT -0.040 -0.020 0.040 0.020 ;
 LAYER M2 ;
 RECT -0.070 -0.020 0.070 0.020 ;
 LAYER C1 ;
 RECT -0.062 -0.042 0.062 0.042 ;
 END VIA02_BAR_H_0_30_22_22_AY_R
 
 VIA VIA02_20_20_20_20_HV_2CUT_H_AY_R DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.105 -0.040 0.105 0.040 ;
 LAYER C1 ;
 RECT -0.105 -0.040 0.105 0.040 ;
 END VIA02_20_20_20_20_HV_2CUT_H_AY_R
 
 VIA VIA02_20_20_20_20_HV_2CUT_V_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.085 0.020 -0.045 ;
 RECT -0.020 0.045 0.020 0.085 ;
 LAYER M2 ;
 RECT -0.040 -0.105 0.040 0.105 ;
 LAYER C1 ;
 RECT -0.040 -0.105 0.040 0.105 ;
 END VIA02_20_20_20_20_HV_2CUT_V_AY_R
 
 VIA VIA02_20_20_30_10_HV_2CUT_H_AY DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.105 -0.040 0.105 0.040 ;
 LAYER C1 ;
 RECT -0.115 -0.030 0.115 0.030 ;
 END VIA02_20_20_30_10_HV_2CUT_H_AY
 
 VIA VIA02_20_20_30_10_HV_2CUT_V_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.085 0.020 -0.045 ;
 RECT -0.020 0.045 0.020 0.085 ;
 LAYER M2 ;
 RECT -0.040 -0.105 0.040 0.105 ;
 LAYER C1 ;
 RECT -0.050 -0.095 0.050 0.095 ;
 END VIA02_20_20_30_10_HV_2CUT_V_AY
 
 VIA VIA02_20_20_30_30_HV_2CUT_H_AY_R DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.105 -0.040 0.105 0.040 ;
 LAYER C1 ;
 RECT -0.115 -0.050 0.115 0.050 ;
 END VIA02_20_20_30_30_HV_2CUT_H_AY_R
 
 VIA VIA02_20_20_30_30_HV_2CUT_V_AY_R DEFAULT
 LAYER AY ;
 RECT -0.020 -0.085 0.020 -0.045 ;
 RECT -0.020 0.045 0.020 0.085 ;
 LAYER M2 ;
 RECT -0.040 -0.105 0.040 0.105 ;
 LAYER C1 ;
 RECT -0.050 -0.115 0.050 0.115 ;
 END VIA02_20_20_30_30_HV_2CUT_V_AY_R
 
 VIA VIA02_0_30_20_20_HV_2CUT_H_AY DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.020 0.115 0.020 ;
 LAYER C1 ;
 RECT -0.105 -0.040 0.105 0.040 ;
 END VIA02_0_30_20_20_HV_2CUT_H_AY
 
 VIA VIA02_0_30_30_10_HV_2CUT_H_AY DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.020 0.115 0.020 ;
 LAYER C1 ;
 RECT -0.115 -0.030 0.115 0.030 ;
 END VIA02_0_30_30_10_HV_2CUT_H_AY
 
 VIA VIA02_0_30_30_30_HV_2CUT_H_AY DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.020 0.115 0.020 ;
 LAYER C1 ;
 RECT -0.115 -0.050 0.115 0.050 ;
 END VIA02_0_30_30_30_HV_2CUT_H_AY
 
 VIA VIA02_10_30_20_20_HV_2CUT_H_AY DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.030 0.115 0.030 ;
 LAYER C1 ;
 RECT -0.105 -0.040 0.105 0.040 ;
 END VIA02_10_30_20_20_HV_2CUT_H_AY
 
 VIA VIA02_10_30_20_20_HV_2CUT_V_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.085 0.020 -0.045 ;
 RECT -0.020 0.045 0.020 0.085 ;
 LAYER M2 ;
 RECT -0.050 -0.095 0.050 0.095 ;
 LAYER C1 ;
 RECT -0.040 -0.105 0.040 0.105 ;
 END VIA02_10_30_20_20_HV_2CUT_V_AY
 
 VIA VIA02_10_30_30_10_HV_2CUT_H_AY DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.030 0.115 0.030 ;
 LAYER C1 ;
 RECT -0.115 -0.030 0.115 0.030 ;
 END VIA02_10_30_30_10_HV_2CUT_H_AY
 
 VIA VIA02_10_30_30_10_HV_2CUT_V_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.085 0.020 -0.045 ;
 RECT -0.020 0.045 0.020 0.085 ;
 LAYER M2 ;
 RECT -0.050 -0.095 0.050 0.095 ;
 LAYER C1 ;
 RECT -0.050 -0.095 0.050 0.095 ;
 END VIA02_10_30_30_10_HV_2CUT_V_AY
 
 VIA VIA02_10_30_30_30_HV_2CUT_H_AY DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.030 0.115 0.030 ;
 LAYER C1 ;
 RECT -0.115 -0.050 0.115 0.050 ;
 END VIA02_10_30_30_30_HV_2CUT_H_AY
 
 VIA VIA02_10_30_30_30_HV_2CUT_V_AY DEFAULT
 LAYER AY ;
 RECT -0.020 -0.085 0.020 -0.045 ;
 RECT -0.020 0.045 0.020 0.085 ;
 LAYER M2 ;
 RECT -0.050 -0.095 0.050 0.095 ;
 LAYER C1 ;
 RECT -0.050 -0.115 0.050 0.115 ;
 END VIA02_10_30_30_30_HV_2CUT_V_AY
 
 VIA VIA02_0_30_2_34_HV_2CUT_H_AY_R DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.020 0.115 0.020 ;
 LAYER C1 ;
 RECT -0.087 -0.054 0.087 0.054 ;
 END VIA02_0_30_2_34_HV_2CUT_H_AY_R
 
 VIA VIA02_0_30_2_53_HV_2CUT_H_AY_R DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.020 0.115 0.020 ;
 LAYER C1 ;
 RECT -0.087 -0.073 0.087 0.073 ;
 END VIA02_0_30_2_53_HV_2CUT_H_AY_R
 
 VIA VIA02_0_30_2_63_HV_2CUT_H_AY_R DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.020 0.115 0.020 ;
 LAYER C1 ;
 RECT -0.087 -0.083 0.087 0.083 ;
 END VIA02_0_30_2_63_HV_2CUT_H_AY_R
 
 VIA VIA02_0_30_7_30_HV_2CUT_H_AY_R DEFAULT
 LAYER AY ;
 RECT -0.085 -0.020 -0.045 0.020 ;
 RECT 0.045 -0.020 0.085 0.020 ;
 LAYER M2 ;
 RECT -0.115 -0.020 0.115 0.020 ;
 LAYER C1 ;
 RECT -0.092 -0.050 0.092 0.050 ;
 END VIA02_0_30_7_30_HV_2CUT_H_AY_R
 
 VIA VIA02_20_20_20_20_XX_4CUT_AY DEFAULT
 LAYER AY ;
 RECT -0.085 -0.085 -0.045 -0.045 ;
 RECT 0.045 -0.085 0.085 -0.045 ;
 RECT -0.085 0.045 -0.045 0.085 ;
 RECT 0.045 0.045 0.085 0.085 ;
 LAYER M2 ;
 RECT -0.105 -0.105 0.105 0.105 ;
 LAYER C1 ;
 RECT -0.105 -0.105 0.105 0.105 ;
 END VIA02_20_20_20_20_XX_4CUT_AY
 
VIARULE VIA02_GEN_0_30_2_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.000 ;
  LAYER C1 ;
    ENCLOSURE 0.002 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_0_30_2_35_HV_AY 

VIARULE VIA02_GEN_0_30_3_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.000 ;
  LAYER C1 ;
    ENCLOSURE 0.003 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_0_30_3_35_HV_AY 

VIARULE VIA02_GEN_0_30_5_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.000 ;
  LAYER C1 ;
    ENCLOSURE 0.005 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_0_30_5_35_HV_AY 

VIARULE VIA02_GEN_0_30_7_30_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.000 ;
  LAYER C1 ;
    ENCLOSURE 0.007 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_0_30_7_30_HV_AY 

VIARULE VIA02_GEN_0_30_10_30_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.000 ;
  LAYER C1 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_0_30_10_30_HV_AY 

VIARULE VIA02_GEN_3_30_2_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.003 ;
  LAYER C1 ;
    ENCLOSURE 0.002 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_3_30_2_35_HV_AY 

VIARULE VIA02_GEN_3_30_3_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.003 ;
  LAYER C1 ;
    ENCLOSURE 0.003 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_3_30_3_35_HV_AY 

VIARULE VIA02_GEN_3_30_5_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.003 ;
  LAYER C1 ;
    ENCLOSURE 0.005 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_3_30_5_35_HV_AY 

VIARULE VIA02_GEN_3_30_7_30_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.003 ;
  LAYER C1 ;
    ENCLOSURE 0.007 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_3_30_7_30_HV_AY 

VIARULE VIA02_GEN_3_30_10_30_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.003 ;
  LAYER C1 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_3_30_10_30_HV_AY 

VIARULE VIA02_GEN_5_30_2_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER C1 ;
    ENCLOSURE 0.002 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_5_30_2_35_HV_AY 

VIARULE VIA02_GEN_5_30_3_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER C1 ;
    ENCLOSURE 0.003 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_5_30_3_35_HV_AY 

VIARULE VIA02_GEN_5_30_5_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER C1 ;
    ENCLOSURE 0.005 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_5_30_5_35_HV_AY 

VIARULE VIA02_GEN_5_30_7_30_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER C1 ;
    ENCLOSURE 0.007 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_5_30_7_30_HV_AY 

VIARULE VIA02_GEN_5_30_10_30_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER C1 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_5_30_10_30_HV_AY 

VIARULE VIA02_GEN_10_25_2_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C1 ;
    ENCLOSURE 0.002 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_10_25_2_35_HV_AY 

VIARULE VIA02_GEN_10_25_3_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C1 ;
    ENCLOSURE 0.003 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_10_25_3_35_HV_AY 

VIARULE VIA02_GEN_10_25_5_35_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C1 ;
    ENCLOSURE 0.005 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_10_25_5_35_HV_AY 

VIARULE VIA02_GEN_10_25_7_30_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C1 ;
    ENCLOSURE 0.007 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_10_25_7_30_HV_AY 

VIARULE VIA02_GEN_10_25_10_30_HV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C1 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_10_25_10_30_HV_AY 

VIARULE VIA02_GEN_20_20_2_35_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C1 ;
    ENCLOSURE 0.002 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_20_20_2_35_XV_AY 

VIARULE VIA02_GEN_20_20_3_35_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C1 ;
    ENCLOSURE 0.003 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_20_20_3_35_XV_AY 

VIARULE VIA02_GEN_20_20_5_35_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C1 ;
    ENCLOSURE 0.005 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_20_20_5_35_XV_AY 

VIARULE VIA02_GEN_20_20_7_30_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C1 ;
    ENCLOSURE 0.007 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_20_20_7_30_XV_AY 

VIARULE VIA02_GEN_20_20_10_30_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C1 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_20_20_10_30_XV_AY 

VIARULE VIA02_GEN_30_30_2_35_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.030 ;
  LAYER C1 ;
    ENCLOSURE 0.002 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_30_30_2_35_XV_AY 

VIARULE VIA02_GEN_30_30_3_35_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.030 ;
  LAYER C1 ;
    ENCLOSURE 0.003 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_30_30_3_35_XV_AY 

VIARULE VIA02_GEN_30_30_5_35_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.030 ;
  LAYER C1 ;
    ENCLOSURE 0.005 0.035 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_30_30_5_35_XV_AY 

VIARULE VIA02_GEN_30_30_7_30_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.030 ;
  LAYER C1 ;
    ENCLOSURE 0.007 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_30_30_7_30_XV_AY 

VIARULE VIA02_GEN_30_30_10_30_XV_AY GENERATE
  LAYER M2 ;
    ENCLOSURE 0.030 0.030 ;
  LAYER C1 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER AY ;
    RECT -0.020 -0.020 0.020 0.020 ;
    SPACING 0.130 BY 0.130 ;
END  VIA02_GEN_30_30_10_30_XV_AY 

#------------------------------------------------------------
#  A1 VIA SECTION 
#------------------------------------------------------------
 VIA VIA03 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA03
 
 VIA VIA03_0_25_0_32_VV_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA03_0_25_0_32_VV_A1
 
 VIA VIA03_0_25_4_20_VH_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA03_0_25_4_20_VH_A1
 
 VIA VIA03_0_25_4_20_VV_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA03_0_25_4_20_VV_A1
 
 VIA VIA03_0_25_18_18_VX_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA03_0_25_18_18_VX_A1
 
 VIA VIA03_4_20_0_32_VH_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA03_4_20_0_32_VH_A1
 
 VIA VIA03_4_20_0_32_VV_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA03_4_20_0_32_VV_A1
 
 VIA VIA03_4_20_4_20_VH_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA03_4_20_4_20_VH_A1
 
 VIA VIA03_4_20_4_20_VV_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA03_4_20_4_20_VV_A1
 
 VIA VIA03_4_20_18_18_VX_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA03_4_20_18_18_VX_A1
 
 VIA VIA03_BAR_V_0_36_23_23_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C1 ;
 RECT -0.022 -0.081 0.022 0.081 ;
 LAYER C2 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA03_BAR_V_0_36_23_23_A1
 
 VIA VIA03_BAR_V_9_27_23_23_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C1 ;
 RECT -0.031 -0.072 0.031 0.072 ;
 LAYER C2 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA03_BAR_V_9_27_23_23_A1
 
 VIA VIA03_BAR_V_18_18_23_23_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C1 ;
 RECT -0.040 -0.063 0.040 0.063 ;
 LAYER C2 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA03_BAR_V_18_18_23_23_A1
 
 VIA VIA03_BAR_H_23_23_0_36_A1 DEFAULT
 LAYER A1 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C1 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C2 ;
 RECT -0.081 -0.022 0.081 0.022 ;
 END VIA03_BAR_H_23_23_0_36_A1
 
 VIA VIA03_BAR_H_23_23_9_27_A1 DEFAULT
 LAYER A1 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C1 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C2 ;
 RECT -0.072 -0.031 0.072 0.031 ;
 END VIA03_BAR_H_23_23_9_27_A1
 
 VIA VIA03_BAR_H_23_23_18_18_A1 DEFAULT
 LAYER A1 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C1 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C2 ;
 RECT -0.063 -0.040 0.063 0.040 ;
 END VIA03_BAR_H_23_23_18_18_A1
 
 VIA VIA03_BAR_H_23_23_23_23_A1 DEFAULT
 LAYER A1 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C1 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C2 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA03_BAR_H_23_23_23_23_A1
 
 VIA VIA03_BAR_V_23_23_23_23_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C1 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C2 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA03_BAR_V_23_23_23_23_A1
 
 VIA VIA03_0_25_0_53_VH_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA03_0_25_0_53_VH_A1_R
 
 VIA VIA03_0_25_0_53_VV_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA03_0_25_0_53_VV_A1_R
 
 VIA VIA03_0_25_0_63_VH_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA03_0_25_0_63_VH_A1_R
 
 VIA VIA03_0_25_0_63_VV_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C2 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA03_0_25_0_63_VV_A1_R
 
 VIA VIA03_4_20_0_53_VH_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA03_4_20_0_53_VH_A1_R
 
 VIA VIA03_4_20_0_53_VV_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA03_4_20_0_53_VV_A1_R
 
 VIA VIA03_4_20_0_63_VH_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA03_4_20_0_63_VH_A1_R
 
 VIA VIA03_4_20_0_63_VV_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C1 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C2 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA03_4_20_0_63_VV_A1_R
 
 VIA VIA03_BAR_H_9_27_0_47_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C1 ;
 RECT -0.072 -0.031 0.072 0.031 ;
 LAYER C2 ;
 RECT -0.092 -0.022 0.092 0.022 ;
 END VIA03_BAR_H_9_27_0_47_A1_R
 
 VIA VIA03_BAR_H_18_18_0_47_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C1 ;
 RECT -0.063 -0.040 0.063 0.040 ;
 LAYER C2 ;
 RECT -0.092 -0.022 0.092 0.022 ;
 END VIA03_BAR_H_18_18_0_47_A1_R
 
 VIA VIA03_BAR_V_0_36_22_22_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C1 ;
 RECT -0.022 -0.081 0.022 0.081 ;
 LAYER C2 ;
 RECT -0.044 -0.067 0.044 0.067 ;
 END VIA03_BAR_V_0_36_22_22_A1_R
 
 VIA VIA03_0_25_0_32_VH_2CUT_H_A1 DEFAULT
 LAYER A1 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C1 ;
 RECT -0.085 -0.047 0.085 0.047 ;
 LAYER C2 ;
 RECT -0.117 -0.022 0.117 0.022 ;
 END VIA03_0_25_0_32_VH_2CUT_H_A1
 
 VIA VIA03_0_25_4_20_VH_2CUT_V_A1 DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C1 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C2 ;
 RECT -0.042 -0.089 0.042 0.089 ;
 END VIA03_0_25_4_20_VH_2CUT_V_A1
 
 VIA VIA03_0_25_18_18_VH_2CUT_V_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C1 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C2 ;
 RECT -0.040 -0.103 0.040 0.103 ;
 END VIA03_0_25_18_18_VH_2CUT_V_A1_R
 
 VIA VIA03_0_25_0_32_VH_2CUT_V_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C1 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C2 ;
 RECT -0.054 -0.085 0.054 0.085 ;
 END VIA03_0_25_0_32_VH_2CUT_V_A1_R
 
 VIA VIA03_0_25_0_53_VH_2CUT_V_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C1 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C2 ;
 RECT -0.075 -0.085 0.075 0.085 ;
 END VIA03_0_25_0_53_VH_2CUT_V_A1_R
 
 VIA VIA03_0_25_0_63_VX_2CUT_V_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C1 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C2 ;
 RECT -0.085 -0.085 0.085 0.085 ;
 END VIA03_0_25_0_63_VX_2CUT_V_A1_R
 
 VIA VIA03_0_25_10_20_VH_2CUT_V_A1_R DEFAULT
 LAYER A1 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C1 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C2 ;
 RECT -0.042 -0.095 0.042 0.095 ;
 END VIA03_0_25_10_20_VH_2CUT_V_A1_R
 
 VIA VIA03_0_25_10_20_VH_4CUT_A1 DEFAULT
 LAYER A1 ;
 RECT -0.085 -0.085 -0.041 -0.041 ;
 RECT 0.041 -0.085 0.085 -0.041 ;
 RECT -0.085 0.041 -0.041 0.085 ;
 RECT 0.041 0.041 0.085 0.085 ;
 LAYER C1 ;
 RECT -0.085 -0.110 0.085 0.110 ;
 LAYER C2 ;
 RECT -0.105 -0.095 0.105 0.095 ;
 END VIA03_0_25_10_20_VH_4CUT_A1
 
VIARULE VIA03_GEN_0_25_0_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_0_25_0_32_VH_A1 

VIARULE VIA03_GEN_0_25_2_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_0_25_2_32_VH_A1 

VIARULE VIA03_GEN_0_25_5_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_0_25_5_30_VH_A1 

VIARULE VIA03_GEN_0_25_10_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_0_25_10_30_VH_A1 

VIARULE VIA03_GEN_0_25_15_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_0_25_15_30_VH_A1 

VIARULE VIA03_GEN_0_25_20_20_VX_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_0_25_20_20_VX_A1 

VIARULE VIA03_GEN_0_25_20_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_0_25_20_30_VH_A1 

VIARULE VIA03_GEN_2_25_0_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_2_25_0_32_VH_A1 

VIARULE VIA03_GEN_2_25_2_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_2_25_2_32_VH_A1 

VIARULE VIA03_GEN_2_25_5_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_2_25_5_30_VH_A1 

VIARULE VIA03_GEN_2_25_10_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_2_25_10_30_VH_A1 

VIARULE VIA03_GEN_2_25_15_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_2_25_15_30_VH_A1 

VIARULE VIA03_GEN_2_25_20_20_VX_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_2_25_20_20_VX_A1 

VIARULE VIA03_GEN_2_25_20_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_2_25_20_30_VH_A1 

VIARULE VIA03_GEN_5_25_0_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_5_25_0_32_VH_A1 

VIARULE VIA03_GEN_5_25_2_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_5_25_2_32_VH_A1 

VIARULE VIA03_GEN_5_25_5_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_5_25_5_30_VH_A1 

VIARULE VIA03_GEN_5_25_10_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_5_25_10_30_VH_A1 

VIARULE VIA03_GEN_5_25_15_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_5_25_15_30_VH_A1 

VIARULE VIA03_GEN_5_25_20_20_VX_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_5_25_20_20_VX_A1 

VIARULE VIA03_GEN_5_25_20_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_5_25_20_30_VH_A1 

VIARULE VIA03_GEN_10_25_0_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_10_25_0_32_VH_A1 

VIARULE VIA03_GEN_10_25_2_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_10_25_2_32_VH_A1 

VIARULE VIA03_GEN_10_25_5_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_10_25_5_30_VH_A1 

VIARULE VIA03_GEN_10_25_10_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_10_25_10_30_VH_A1 

VIARULE VIA03_GEN_10_25_15_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_10_25_15_30_VH_A1 

VIARULE VIA03_GEN_10_25_20_20_VX_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_10_25_20_20_VX_A1 

VIARULE VIA03_GEN_10_25_20_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_10_25_20_30_VH_A1 

VIARULE VIA03_GEN_15_25_0_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_15_25_0_32_VH_A1 

VIARULE VIA03_GEN_15_25_2_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_15_25_2_32_VH_A1 

VIARULE VIA03_GEN_15_25_5_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_15_25_5_30_VH_A1 

VIARULE VIA03_GEN_15_25_10_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_15_25_10_30_VH_A1 

VIARULE VIA03_GEN_15_25_15_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_15_25_15_30_VH_A1 

VIARULE VIA03_GEN_15_25_20_20_VX_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_15_25_20_20_VX_A1 

VIARULE VIA03_GEN_15_25_20_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_15_25_20_30_VH_A1 

VIARULE VIA03_GEN_20_30_0_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_20_30_0_32_VH_A1 

VIARULE VIA03_GEN_20_30_2_32_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C2 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_20_30_2_32_VH_A1 

VIARULE VIA03_GEN_20_30_5_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_20_30_5_30_VH_A1 

VIARULE VIA03_GEN_20_30_10_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_20_30_10_30_VH_A1 

VIARULE VIA03_GEN_20_30_15_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_20_30_15_30_VH_A1 

VIARULE VIA03_GEN_20_30_20_20_VX_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_20_30_20_20_VX_A1 

VIARULE VIA03_GEN_20_30_20_30_VH_A1 GENERATE
  LAYER C1 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A1 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA03_GEN_20_30_20_30_VH_A1 

#------------------------------------------------------------
#  A2 VIA SECTION 
#------------------------------------------------------------
 VIA VIA04_0_25_0_32_HH_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA04_0_25_0_32_HH_A2
 
 VIA VIA04 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA04
 
 VIA VIA04_0_25_4_20_HH_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA04_0_25_4_20_HH_A2
 
 VIA VIA04_0_25_4_20_HV_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA04_0_25_4_20_HV_A2
 
 VIA VIA04_0_25_18_18_HX_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA04_0_25_18_18_HX_A2
 
 VIA VIA04_4_20_0_32_HH_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA04_4_20_0_32_HH_A2
 
 VIA VIA04_4_20_0_32_HV_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA04_4_20_0_32_HV_A2
 
 VIA VIA04_4_20_4_20_HH_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA04_4_20_4_20_HH_A2
 
 VIA VIA04_4_20_4_20_HV_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA04_4_20_4_20_HV_A2
 
 VIA VIA04_4_20_18_18_HX_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA04_4_20_18_18_HX_A2
 
 VIA VIA04_18_18_0_32_XH_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA04_18_18_0_32_XH_A2
 
 VIA VIA04_18_18_0_32_XV_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA04_18_18_0_32_XV_A2
 
 VIA VIA04_18_18_4_20_XH_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA04_18_18_4_20_XH_A2
 
 VIA VIA04_18_18_4_20_XV_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA04_18_18_4_20_XV_A2
 
 VIA VIA04_18_18_18_18_XX_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA04_18_18_18_18_XX_A2
 
 VIA VIA04_BAR_H_0_36_23_23_A2 DEFAULT
 LAYER A2 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C2 ;
 RECT -0.081 -0.022 0.081 0.022 ;
 LAYER C3 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA04_BAR_H_0_36_23_23_A2
 
 VIA VIA04_BAR_H_9_27_23_23_A2 DEFAULT
 LAYER A2 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C2 ;
 RECT -0.072 -0.031 0.072 0.031 ;
 LAYER C3 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA04_BAR_H_9_27_23_23_A2
 
 VIA VIA04_BAR_H_18_18_23_23_A2 DEFAULT
 LAYER A2 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C2 ;
 RECT -0.063 -0.040 0.063 0.040 ;
 LAYER C3 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA04_BAR_H_18_18_23_23_A2
 
 VIA VIA04_BAR_V_23_23_0_36_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C2 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C3 ;
 RECT -0.022 -0.081 0.022 0.081 ;
 END VIA04_BAR_V_23_23_0_36_A2
 
 VIA VIA04_BAR_V_23_23_9_27_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C2 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C3 ;
 RECT -0.031 -0.072 0.031 0.072 ;
 END VIA04_BAR_V_23_23_9_27_A2
 
 VIA VIA04_BAR_V_23_23_18_18_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C2 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C3 ;
 RECT -0.040 -0.063 0.040 0.063 ;
 END VIA04_BAR_V_23_23_18_18_A2
 
 VIA VIA04_BAR_H_23_23_23_23_A2 DEFAULT
 LAYER A2 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C2 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C3 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA04_BAR_H_23_23_23_23_A2
 
 VIA VIA04_BAR_V_23_23_23_23_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C2 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C3 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA04_BAR_V_23_23_23_23_A2
 
 VIA VIA04_0_25_0_53_HH_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA04_0_25_0_53_HH_A2_R
 
 VIA VIA04_0_25_0_53_HV_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA04_0_25_0_53_HV_A2_R
 
 VIA VIA04_0_25_0_63_HH_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA04_0_25_0_63_HH_A2_R
 
 VIA VIA04_0_25_0_63_HV_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA04_0_25_0_63_HV_A2_R
 
 VIA VIA04_4_20_0_53_HH_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA04_4_20_0_53_HH_A2_R
 
 VIA VIA04_4_20_0_53_HV_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA04_4_20_0_53_HV_A2_R
 
 VIA VIA04_4_20_0_63_HH_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA04_4_20_0_63_HH_A2_R
 
 VIA VIA04_4_20_0_63_HV_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C3 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA04_4_20_0_63_HV_A2_R
 
 VIA VIA04_18_18_0_53_XH_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA04_18_18_0_53_XH_A2_R
 
 VIA VIA04_18_18_0_53_XV_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA04_18_18_0_53_XV_A2_R
 
 VIA VIA04_18_18_0_63_XH_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA04_18_18_0_63_XH_A2_R
 
 VIA VIA04_18_18_0_63_XV_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C2 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C3 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA04_18_18_0_63_XV_A2_R
 
 VIA VIA04_BAR_V_9_27_0_47_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C2 ;
 RECT -0.031 -0.072 0.031 0.072 ;
 LAYER C3 ;
 RECT -0.022 -0.092 0.022 0.092 ;
 END VIA04_BAR_V_9_27_0_47_A2_R
 
 VIA VIA04_BAR_V_18_18_0_47_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C2 ;
 RECT -0.040 -0.063 0.040 0.063 ;
 LAYER C3 ;
 RECT -0.022 -0.092 0.022 0.092 ;
 END VIA04_BAR_V_18_18_0_47_A2_R
 
 VIA VIA04_BAR_H_0_36_22_22_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C2 ;
 RECT -0.081 -0.022 0.081 0.022 ;
 LAYER C3 ;
 RECT -0.067 -0.044 0.067 0.044 ;
 END VIA04_BAR_H_0_36_22_22_A2_R
 
 VIA VIA04_0_25_0_32_HV_2CUT_V_A2 DEFAULT
 LAYER A2 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C2 ;
 RECT -0.047 -0.085 0.047 0.085 ;
 LAYER C3 ;
 RECT -0.022 -0.117 0.022 0.117 ;
 END VIA04_0_25_0_32_HV_2CUT_V_A2
 
 VIA VIA04_0_25_4_20_HV_2CUT_H_A2 DEFAULT
 LAYER A2 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C2 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C3 ;
 RECT -0.089 -0.042 0.089 0.042 ;
 END VIA04_0_25_4_20_HV_2CUT_H_A2
 
 VIA VIA04_0_25_18_18_HV_2CUT_H_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C2 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C3 ;
 RECT -0.103 -0.040 0.103 0.040 ;
 END VIA04_0_25_18_18_HV_2CUT_H_A2_R
 
 VIA VIA04_0_25_0_32_HV_2CUT_H_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C2 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C3 ;
 RECT -0.085 -0.054 0.085 0.054 ;
 END VIA04_0_25_0_32_HV_2CUT_H_A2_R
 
 VIA VIA04_0_25_0_53_HV_2CUT_H_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C2 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C3 ;
 RECT -0.085 -0.075 0.085 0.075 ;
 END VIA04_0_25_0_53_HV_2CUT_H_A2_R
 
 VIA VIA04_0_25_0_63_HX_2CUT_H_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C2 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C3 ;
 RECT -0.085 -0.085 0.085 0.085 ;
 END VIA04_0_25_0_63_HX_2CUT_H_A2_R
 
 VIA VIA04_0_25_10_20_HV_2CUT_H_A2_R DEFAULT
 LAYER A2 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C2 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C3 ;
 RECT -0.095 -0.042 0.095 0.042 ;
 END VIA04_0_25_10_20_HV_2CUT_H_A2_R
 
 VIA VIA04_0_25_10_20_HV_4CUT_A2 DEFAULT
 LAYER A2 ;
 RECT -0.085 -0.085 -0.041 -0.041 ;
 RECT 0.041 -0.085 0.085 -0.041 ;
 RECT -0.085 0.041 -0.041 0.085 ;
 RECT 0.041 0.041 0.085 0.085 ;
 LAYER C2 ;
 RECT -0.110 -0.085 0.110 0.085 ;
 LAYER C3 ;
 RECT -0.095 -0.105 0.095 0.105 ;
 END VIA04_0_25_10_20_HV_4CUT_A2
 
VIARULE VIA04_GEN_0_25_0_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C3 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_0_25_0_32_HV_A2 

VIARULE VIA04_GEN_0_25_2_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C3 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_0_25_2_32_HV_A2 

VIARULE VIA04_GEN_0_25_5_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C3 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_0_25_5_30_HV_A2 

VIARULE VIA04_GEN_0_25_10_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C3 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_0_25_10_30_HV_A2 

VIARULE VIA04_GEN_0_25_15_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C3 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_0_25_15_30_HV_A2 

VIARULE VIA04_GEN_0_25_20_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_0_25_20_30_HV_A2 

VIARULE VIA04_GEN_2_25_0_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C3 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_2_25_0_32_HV_A2 

VIARULE VIA04_GEN_2_25_2_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C3 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_2_25_2_32_HV_A2 

VIARULE VIA04_GEN_2_25_5_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C3 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_2_25_5_30_HV_A2 

VIARULE VIA04_GEN_2_25_10_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C3 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_2_25_10_30_HV_A2 

VIARULE VIA04_GEN_2_25_15_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C3 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_2_25_15_30_HV_A2 

VIARULE VIA04_GEN_2_25_20_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_2_25_20_30_HV_A2 

VIARULE VIA04_GEN_5_25_0_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C3 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_5_25_0_32_HV_A2 

VIARULE VIA04_GEN_5_25_2_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C3 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_5_25_2_32_HV_A2 

VIARULE VIA04_GEN_5_25_5_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C3 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_5_25_5_30_HV_A2 

VIARULE VIA04_GEN_5_25_10_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C3 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_5_25_10_30_HV_A2 

VIARULE VIA04_GEN_5_25_15_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C3 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_5_25_15_30_HV_A2 

VIARULE VIA04_GEN_5_25_20_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_5_25_20_30_HV_A2 

VIARULE VIA04_GEN_10_25_0_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C3 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_10_25_0_32_HV_A2 

VIARULE VIA04_GEN_10_25_2_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C3 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_10_25_2_32_HV_A2 

VIARULE VIA04_GEN_10_25_5_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C3 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_10_25_5_30_HV_A2 

VIARULE VIA04_GEN_10_25_10_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C3 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_10_25_10_30_HV_A2 

VIARULE VIA04_GEN_10_25_15_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C3 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_10_25_15_30_HV_A2 

VIARULE VIA04_GEN_10_25_20_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_10_25_20_30_HV_A2 

VIARULE VIA04_GEN_15_25_0_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C3 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_15_25_0_32_HV_A2 

VIARULE VIA04_GEN_15_25_2_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C3 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_15_25_2_32_HV_A2 

VIARULE VIA04_GEN_15_25_5_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C3 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_15_25_5_30_HV_A2 

VIARULE VIA04_GEN_15_25_10_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C3 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_15_25_10_30_HV_A2 

VIARULE VIA04_GEN_15_25_15_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C3 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_15_25_15_30_HV_A2 

VIARULE VIA04_GEN_15_25_20_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_15_25_20_30_HV_A2 

VIARULE VIA04_GEN_20_20_0_32_XV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_20_0_32_XV_A2 

VIARULE VIA04_GEN_20_20_2_32_XV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_20_2_32_XV_A2 

VIARULE VIA04_GEN_20_20_5_30_XV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_20_5_30_XV_A2 

VIARULE VIA04_GEN_20_20_10_30_XV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_20_10_30_XV_A2 

VIARULE VIA04_GEN_20_20_15_30_XV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_20_15_30_XV_A2 

VIARULE VIA04_GEN_20_20_20_30_XV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_20_20_30_XV_A2 

VIARULE VIA04_GEN_20_30_0_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_30_0_32_HV_A2 

VIARULE VIA04_GEN_20_30_2_32_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_30_2_32_HV_A2 

VIARULE VIA04_GEN_20_30_5_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_30_5_30_HV_A2 

VIARULE VIA04_GEN_20_30_10_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_30_10_30_HV_A2 

VIARULE VIA04_GEN_20_30_15_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_30_15_30_HV_A2 

VIARULE VIA04_GEN_20_30_20_30_HV_A2 GENERATE
  LAYER C2 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A2 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA04_GEN_20_30_20_30_HV_A2 

#------------------------------------------------------------
#  A3 VIA SECTION 
#------------------------------------------------------------
 VIA VIA05 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA05
 
 VIA VIA05_0_25_0_32_VV_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA05_0_25_0_32_VV_A3
 
 VIA VIA05_0_25_4_20_VH_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA05_0_25_4_20_VH_A3
 
 VIA VIA05_0_25_4_20_VV_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA05_0_25_4_20_VV_A3
 
 VIA VIA05_0_25_18_18_VX_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA05_0_25_18_18_VX_A3
 
 VIA VIA05_4_20_0_32_VH_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA05_4_20_0_32_VH_A3
 
 VIA VIA05_4_20_0_32_VV_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA05_4_20_0_32_VV_A3
 
 VIA VIA05_4_20_4_20_VH_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA05_4_20_4_20_VH_A3
 
 VIA VIA05_4_20_4_20_VV_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA05_4_20_4_20_VV_A3
 
 VIA VIA05_4_20_18_18_VX_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA05_4_20_18_18_VX_A3
 
 VIA VIA05_BAR_V_0_36_23_23_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C3 ;
 RECT -0.022 -0.081 0.022 0.081 ;
 LAYER C4 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA05_BAR_V_0_36_23_23_A3
 
 VIA VIA05_BAR_V_9_27_23_23_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C3 ;
 RECT -0.031 -0.072 0.031 0.072 ;
 LAYER C4 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA05_BAR_V_9_27_23_23_A3
 
 VIA VIA05_BAR_V_18_18_23_23_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C3 ;
 RECT -0.040 -0.063 0.040 0.063 ;
 LAYER C4 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA05_BAR_V_18_18_23_23_A3
 
 VIA VIA05_BAR_H_23_23_0_36_A3 DEFAULT
 LAYER A3 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C3 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C4 ;
 RECT -0.081 -0.022 0.081 0.022 ;
 END VIA05_BAR_H_23_23_0_36_A3
 
 VIA VIA05_BAR_H_23_23_9_27_A3 DEFAULT
 LAYER A3 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C3 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C4 ;
 RECT -0.072 -0.031 0.072 0.031 ;
 END VIA05_BAR_H_23_23_9_27_A3
 
 VIA VIA05_BAR_H_23_23_18_18_A3 DEFAULT
 LAYER A3 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C3 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C4 ;
 RECT -0.063 -0.040 0.063 0.040 ;
 END VIA05_BAR_H_23_23_18_18_A3
 
 VIA VIA05_BAR_H_23_23_23_23_A3 DEFAULT
 LAYER A3 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C3 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C4 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA05_BAR_H_23_23_23_23_A3
 
 VIA VIA05_BAR_V_23_23_23_23_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C3 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C4 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA05_BAR_V_23_23_23_23_A3
 
 VIA VIA05_0_25_0_53_VH_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA05_0_25_0_53_VH_A3_R
 
 VIA VIA05_0_25_0_53_VV_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA05_0_25_0_53_VV_A3_R
 
 VIA VIA05_0_25_0_63_VH_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA05_0_25_0_63_VH_A3_R
 
 VIA VIA05_0_25_0_63_VV_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.022 -0.047 0.022 0.047 ;
 LAYER C4 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA05_0_25_0_63_VV_A3_R
 
 VIA VIA05_4_20_0_53_VH_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA05_4_20_0_53_VH_A3_R
 
 VIA VIA05_4_20_0_53_VV_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA05_4_20_0_53_VV_A3_R
 
 VIA VIA05_4_20_0_63_VH_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA05_4_20_0_63_VH_A3_R
 
 VIA VIA05_4_20_0_63_VV_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C3 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 LAYER C4 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA05_4_20_0_63_VV_A3_R
 
 VIA VIA05_BAR_H_9_27_0_47_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C3 ;
 RECT -0.072 -0.031 0.072 0.031 ;
 LAYER C4 ;
 RECT -0.092 -0.022 0.092 0.022 ;
 END VIA05_BAR_H_9_27_0_47_A3_R
 
 VIA VIA05_BAR_H_18_18_0_47_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C3 ;
 RECT -0.063 -0.040 0.063 0.040 ;
 LAYER C4 ;
 RECT -0.092 -0.022 0.092 0.022 ;
 END VIA05_BAR_H_18_18_0_47_A3_R
 
 VIA VIA05_BAR_V_0_36_22_22_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C3 ;
 RECT -0.022 -0.081 0.022 0.081 ;
 LAYER C4 ;
 RECT -0.044 -0.067 0.044 0.067 ;
 END VIA05_BAR_V_0_36_22_22_A3_R
 
 VIA VIA05_0_25_0_32_VH_2CUT_H_A3 DEFAULT
 LAYER A3 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C3 ;
 RECT -0.085 -0.047 0.085 0.047 ;
 LAYER C4 ;
 RECT -0.117 -0.022 0.117 0.022 ;
 END VIA05_0_25_0_32_VH_2CUT_H_A3
 
 VIA VIA05_0_25_4_20_VH_2CUT_V_A3 DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C3 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C4 ;
 RECT -0.042 -0.089 0.042 0.089 ;
 END VIA05_0_25_4_20_VH_2CUT_V_A3
 
 VIA VIA05_0_25_18_18_VH_2CUT_V_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C3 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C4 ;
 RECT -0.040 -0.103 0.040 0.103 ;
 END VIA05_0_25_18_18_VH_2CUT_V_A3_R
 
 VIA VIA05_0_25_0_32_VH_2CUT_V_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C3 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C4 ;
 RECT -0.054 -0.085 0.054 0.085 ;
 END VIA05_0_25_0_32_VH_2CUT_V_A3_R
 
 VIA VIA05_0_25_0_53_VH_2CUT_V_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C3 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C4 ;
 RECT -0.075 -0.085 0.075 0.085 ;
 END VIA05_0_25_0_53_VH_2CUT_V_A3_R
 
 VIA VIA05_0_25_0_63_VX_2CUT_V_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C3 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C4 ;
 RECT -0.085 -0.085 0.085 0.085 ;
 END VIA05_0_25_0_63_VX_2CUT_V_A3_R
 
 VIA VIA05_0_25_10_20_VH_2CUT_V_A3_R DEFAULT
 LAYER A3 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C3 ;
 RECT -0.022 -0.110 0.022 0.110 ;
 LAYER C4 ;
 RECT -0.042 -0.095 0.042 0.095 ;
 END VIA05_0_25_10_20_VH_2CUT_V_A3_R
 
 VIA VIA05_0_25_10_20_VH_4CUT_A3 DEFAULT
 LAYER A3 ;
 RECT -0.085 -0.085 -0.041 -0.041 ;
 RECT 0.041 -0.085 0.085 -0.041 ;
 RECT -0.085 0.041 -0.041 0.085 ;
 RECT 0.041 0.041 0.085 0.085 ;
 LAYER C3 ;
 RECT -0.085 -0.110 0.085 0.110 ;
 LAYER C4 ;
 RECT -0.105 -0.095 0.105 0.095 ;
 END VIA05_0_25_10_20_VH_4CUT_A3
 
VIARULE VIA05_GEN_0_25_0_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_0_25_0_32_VH_A3 

VIARULE VIA05_GEN_0_25_2_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_0_25_2_32_VH_A3 

VIARULE VIA05_GEN_0_25_5_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_0_25_5_30_VH_A3 

VIARULE VIA05_GEN_0_25_10_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_0_25_10_30_VH_A3 

VIARULE VIA05_GEN_0_25_15_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_0_25_15_30_VH_A3 

VIARULE VIA05_GEN_0_25_20_20_VX_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_0_25_20_20_VX_A3 

VIARULE VIA05_GEN_0_25_20_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.000 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_0_25_20_30_VH_A3 

VIARULE VIA05_GEN_2_25_0_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_2_25_0_32_VH_A3 

VIARULE VIA05_GEN_2_25_2_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_2_25_2_32_VH_A3 

VIARULE VIA05_GEN_2_25_5_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_2_25_5_30_VH_A3 

VIARULE VIA05_GEN_2_25_10_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_2_25_10_30_VH_A3 

VIARULE VIA05_GEN_2_25_15_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_2_25_15_30_VH_A3 

VIARULE VIA05_GEN_2_25_20_20_VX_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_2_25_20_20_VX_A3 

VIARULE VIA05_GEN_2_25_20_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.002 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_2_25_20_30_VH_A3 

VIARULE VIA05_GEN_5_25_0_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_5_25_0_32_VH_A3 

VIARULE VIA05_GEN_5_25_2_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_5_25_2_32_VH_A3 

VIARULE VIA05_GEN_5_25_5_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_5_25_5_30_VH_A3 

VIARULE VIA05_GEN_5_25_10_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_5_25_10_30_VH_A3 

VIARULE VIA05_GEN_5_25_15_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_5_25_15_30_VH_A3 

VIARULE VIA05_GEN_5_25_20_20_VX_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_5_25_20_20_VX_A3 

VIARULE VIA05_GEN_5_25_20_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.005 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_5_25_20_30_VH_A3 

VIARULE VIA05_GEN_10_25_0_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_10_25_0_32_VH_A3 

VIARULE VIA05_GEN_10_25_2_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_10_25_2_32_VH_A3 

VIARULE VIA05_GEN_10_25_5_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_10_25_5_30_VH_A3 

VIARULE VIA05_GEN_10_25_10_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_10_25_10_30_VH_A3 

VIARULE VIA05_GEN_10_25_15_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_10_25_15_30_VH_A3 

VIARULE VIA05_GEN_10_25_20_20_VX_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_10_25_20_20_VX_A3 

VIARULE VIA05_GEN_10_25_20_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.010 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_10_25_20_30_VH_A3 

VIARULE VIA05_GEN_15_25_0_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_15_25_0_32_VH_A3 

VIARULE VIA05_GEN_15_25_2_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_15_25_2_32_VH_A3 

VIARULE VIA05_GEN_15_25_5_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_15_25_5_30_VH_A3 

VIARULE VIA05_GEN_15_25_10_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_15_25_10_30_VH_A3 

VIARULE VIA05_GEN_15_25_15_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_15_25_15_30_VH_A3 

VIARULE VIA05_GEN_15_25_20_20_VX_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_15_25_20_20_VX_A3 

VIARULE VIA05_GEN_15_25_20_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.015 0.025 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_15_25_20_30_VH_A3 

VIARULE VIA05_GEN_20_30_0_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.000 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_20_30_0_32_VH_A3 

VIARULE VIA05_GEN_20_30_2_32_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C4 ;
    ENCLOSURE 0.032 0.002 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_20_30_2_32_VH_A3 

VIARULE VIA05_GEN_20_30_5_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.005 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_20_30_5_30_VH_A3 

VIARULE VIA05_GEN_20_30_10_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.010 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_20_30_10_30_VH_A3 

VIARULE VIA05_GEN_20_30_15_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.015 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_20_30_15_30_VH_A3 

VIARULE VIA05_GEN_20_30_20_20_VX_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_20_30_20_20_VX_A3 

VIARULE VIA05_GEN_20_30_20_30_VH_A3 GENERATE
  LAYER C3 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER A3 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA05_GEN_20_30_20_30_VH_A3 

#------------------------------------------------------------
#  A4 VIA SECTION 
#------------------------------------------------------------
 VIA VIA06_0_25_0_32_HH_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA06_0_25_0_32_HH_A4
 
 VIA VIA06 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA06
 
 VIA VIA06_0_25_4_20_HH_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA06_0_25_4_20_HH_A4
 
 VIA VIA06_0_25_4_20_HV_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA06_0_25_4_20_HV_A4
 
 VIA VIA06_0_25_18_18_HX_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA06_0_25_18_18_HX_A4
 
 VIA VIA06_4_20_0_32_HH_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA06_4_20_0_32_HH_A4
 
 VIA VIA06_4_20_0_32_HV_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA06_4_20_0_32_HV_A4
 
 VIA VIA06_4_20_4_20_HH_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA06_4_20_4_20_HH_A4
 
 VIA VIA06_4_20_4_20_HV_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA06_4_20_4_20_HV_A4
 
 VIA VIA06_4_20_18_18_HX_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA06_4_20_18_18_HX_A4
 
 VIA VIA06_18_18_0_32_XH_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.054 -0.022 0.054 0.022 ;
 END VIA06_18_18_0_32_XH_A4
 
 VIA VIA06_18_18_0_32_XV_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.022 -0.054 0.022 0.054 ;
 END VIA06_18_18_0_32_XV_A4
 
 VIA VIA06_18_18_4_20_XH_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 END VIA06_18_18_4_20_XH_A4
 
 VIA VIA06_18_18_4_20_XV_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.026 -0.042 0.026 0.042 ;
 END VIA06_18_18_4_20_XV_A4
 
 VIA VIA06_18_18_18_18_XX_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 END VIA06_18_18_18_18_XX_A4
 
 VIA VIA06_BAR_H_0_36_23_23_A4 DEFAULT
 LAYER A4 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C4 ;
 RECT -0.081 -0.022 0.081 0.022 ;
 LAYER C5 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA06_BAR_H_0_36_23_23_A4
 
 VIA VIA06_BAR_H_9_27_23_23_A4 DEFAULT
 LAYER A4 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C4 ;
 RECT -0.072 -0.031 0.072 0.031 ;
 LAYER C5 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA06_BAR_H_9_27_23_23_A4
 
 VIA VIA06_BAR_H_18_18_23_23_A4 DEFAULT
 LAYER A4 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C4 ;
 RECT -0.063 -0.040 0.063 0.040 ;
 LAYER C5 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA06_BAR_H_18_18_23_23_A4
 
 VIA VIA06_BAR_V_23_23_0_36_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C4 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C5 ;
 RECT -0.022 -0.081 0.022 0.081 ;
 END VIA06_BAR_V_23_23_0_36_A4
 
 VIA VIA06_BAR_V_23_23_9_27_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C4 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C5 ;
 RECT -0.031 -0.072 0.031 0.072 ;
 END VIA06_BAR_V_23_23_9_27_A4
 
 VIA VIA06_BAR_V_23_23_18_18_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C4 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C5 ;
 RECT -0.040 -0.063 0.040 0.063 ;
 END VIA06_BAR_V_23_23_18_18_A4
 
 VIA VIA06_BAR_H_23_23_23_23_A4 DEFAULT
 LAYER A4 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C4 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 LAYER C5 ;
 RECT -0.068 -0.045 0.068 0.045 ;
 END VIA06_BAR_H_23_23_23_23_A4
 
 VIA VIA06_BAR_V_23_23_23_23_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C4 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 LAYER C5 ;
 RECT -0.045 -0.068 0.045 0.068 ;
 END VIA06_BAR_V_23_23_23_23_A4
 
 VIA VIA06_0_25_0_53_HH_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA06_0_25_0_53_HH_A4_R
 
 VIA VIA06_0_25_0_53_HV_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA06_0_25_0_53_HV_A4_R
 
 VIA VIA06_0_25_0_63_HH_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA06_0_25_0_63_HH_A4_R
 
 VIA VIA06_0_25_0_63_HV_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.047 -0.022 0.047 0.022 ;
 LAYER C5 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA06_0_25_0_63_HV_A4_R
 
 VIA VIA06_4_20_0_53_HH_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA06_4_20_0_53_HH_A4_R
 
 VIA VIA06_4_20_0_53_HV_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA06_4_20_0_53_HV_A4_R
 
 VIA VIA06_4_20_0_63_HH_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA06_4_20_0_63_HH_A4_R
 
 VIA VIA06_4_20_0_63_HV_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.042 -0.026 0.042 0.026 ;
 LAYER C5 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA06_4_20_0_63_HV_A4_R
 
 VIA VIA06_18_18_0_53_XH_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.075 -0.022 0.075 0.022 ;
 END VIA06_18_18_0_53_XH_A4_R
 
 VIA VIA06_18_18_0_53_XV_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.022 -0.075 0.022 0.075 ;
 END VIA06_18_18_0_53_XV_A4_R
 
 VIA VIA06_18_18_0_63_XH_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.085 -0.022 0.085 0.022 ;
 END VIA06_18_18_0_63_XH_A4_R
 
 VIA VIA06_18_18_0_63_XV_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.022 0.022 0.022 ;
 LAYER C4 ;
 RECT -0.040 -0.040 0.040 0.040 ;
 LAYER C5 ;
 RECT -0.022 -0.085 0.022 0.085 ;
 END VIA06_18_18_0_63_XV_A4_R
 
 VIA VIA06_BAR_V_9_27_0_47_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C4 ;
 RECT -0.031 -0.072 0.031 0.072 ;
 LAYER C5 ;
 RECT -0.022 -0.092 0.022 0.092 ;
 END VIA06_BAR_V_9_27_0_47_A4_R
 
 VIA VIA06_BAR_V_18_18_0_47_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.045 0.022 0.045 ;
 LAYER C4 ;
 RECT -0.040 -0.063 0.040 0.063 ;
 LAYER C5 ;
 RECT -0.022 -0.092 0.022 0.092 ;
 END VIA06_BAR_V_18_18_0_47_A4_R
 
 VIA VIA06_BAR_H_0_36_22_22_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.045 -0.022 0.045 0.022 ;
 LAYER C4 ;
 RECT -0.081 -0.022 0.081 0.022 ;
 LAYER C5 ;
 RECT -0.067 -0.044 0.067 0.044 ;
 END VIA06_BAR_H_0_36_22_22_A4_R
 
 VIA VIA06_0_25_0_32_HV_2CUT_V_A4 DEFAULT
 LAYER A4 ;
 RECT -0.022 -0.085 0.022 -0.041 ;
 RECT -0.022 0.041 0.022 0.085 ;
 LAYER C4 ;
 RECT -0.047 -0.085 0.047 0.085 ;
 LAYER C5 ;
 RECT -0.022 -0.117 0.022 0.117 ;
 END VIA06_0_25_0_32_HV_2CUT_V_A4
 
 VIA VIA06_0_25_4_20_HV_2CUT_H_A4 DEFAULT
 LAYER A4 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C4 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C5 ;
 RECT -0.089 -0.042 0.089 0.042 ;
 END VIA06_0_25_4_20_HV_2CUT_H_A4
 
 VIA VIA06_0_25_18_18_HV_2CUT_H_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C4 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C5 ;
 RECT -0.103 -0.040 0.103 0.040 ;
 END VIA06_0_25_18_18_HV_2CUT_H_A4_R
 
 VIA VIA06_0_25_0_32_HV_2CUT_H_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C4 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C5 ;
 RECT -0.085 -0.054 0.085 0.054 ;
 END VIA06_0_25_0_32_HV_2CUT_H_A4_R
 
 VIA VIA06_0_25_0_53_HV_2CUT_H_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C4 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C5 ;
 RECT -0.085 -0.075 0.085 0.075 ;
 END VIA06_0_25_0_53_HV_2CUT_H_A4_R
 
 VIA VIA06_0_25_0_63_HX_2CUT_H_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C4 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C5 ;
 RECT -0.085 -0.085 0.085 0.085 ;
 END VIA06_0_25_0_63_HX_2CUT_H_A4_R
 
 VIA VIA06_0_25_10_20_HV_2CUT_H_A4_R DEFAULT
 LAYER A4 ;
 RECT -0.085 -0.022 -0.041 0.022 ;
 RECT 0.041 -0.022 0.085 0.022 ;
 LAYER C4 ;
 RECT -0.110 -0.022 0.110 0.022 ;
 LAYER C5 ;
 RECT -0.095 -0.042 0.095 0.042 ;
 END VIA06_0_25_10_20_HV_2CUT_H_A4_R
 
 VIA VIA06_0_25_10_20_HV_4CUT_A4 DEFAULT
 LAYER A4 ;
 RECT -0.085 -0.085 -0.041 -0.041 ;
 RECT 0.041 -0.085 0.085 -0.041 ;
 RECT -0.085 0.041 -0.041 0.085 ;
 RECT 0.041 0.041 0.085 0.085 ;
 LAYER C4 ;
 RECT -0.110 -0.085 0.110 0.085 ;
 LAYER C5 ;
 RECT -0.095 -0.105 0.095 0.105 ;
 END VIA06_0_25_10_20_HV_4CUT_A4
 
VIARULE VIA06_GEN_0_25_0_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C5 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_0_25_0_32_HV_A4 

VIARULE VIA06_GEN_0_25_2_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C5 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_0_25_2_32_HV_A4 

VIARULE VIA06_GEN_0_25_5_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C5 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_0_25_5_30_HV_A4 

VIARULE VIA06_GEN_0_25_10_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C5 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_0_25_10_30_HV_A4 

VIARULE VIA06_GEN_0_25_15_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C5 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_0_25_15_30_HV_A4 

VIARULE VIA06_GEN_0_25_20_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.000 ;
  LAYER C5 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_0_25_20_30_HV_A4 

VIARULE VIA06_GEN_2_25_0_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C5 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_2_25_0_32_HV_A4 

VIARULE VIA06_GEN_2_25_2_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C5 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_2_25_2_32_HV_A4 

VIARULE VIA06_GEN_2_25_5_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C5 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_2_25_5_30_HV_A4 

VIARULE VIA06_GEN_2_25_10_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C5 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_2_25_10_30_HV_A4 

VIARULE VIA06_GEN_2_25_15_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C5 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_2_25_15_30_HV_A4 

VIARULE VIA06_GEN_2_25_20_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.002 ;
  LAYER C5 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_2_25_20_30_HV_A4 

VIARULE VIA06_GEN_5_25_0_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C5 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_5_25_0_32_HV_A4 

VIARULE VIA06_GEN_5_25_2_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C5 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_5_25_2_32_HV_A4 

VIARULE VIA06_GEN_5_25_5_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C5 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_5_25_5_30_HV_A4 

VIARULE VIA06_GEN_5_25_10_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C5 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_5_25_10_30_HV_A4 

VIARULE VIA06_GEN_5_25_15_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C5 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_5_25_15_30_HV_A4 

VIARULE VIA06_GEN_5_25_20_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.005 ;
  LAYER C5 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_5_25_20_30_HV_A4 

VIARULE VIA06_GEN_10_25_0_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C5 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_10_25_0_32_HV_A4 

VIARULE VIA06_GEN_10_25_2_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C5 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_10_25_2_32_HV_A4 

VIARULE VIA06_GEN_10_25_5_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C5 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_10_25_5_30_HV_A4 

VIARULE VIA06_GEN_10_25_10_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C5 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_10_25_10_30_HV_A4 

VIARULE VIA06_GEN_10_25_15_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C5 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_10_25_15_30_HV_A4 

VIARULE VIA06_GEN_10_25_20_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.010 ;
  LAYER C5 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_10_25_20_30_HV_A4 

VIARULE VIA06_GEN_15_25_0_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C5 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_15_25_0_32_HV_A4 

VIARULE VIA06_GEN_15_25_2_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C5 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_15_25_2_32_HV_A4 

VIARULE VIA06_GEN_15_25_5_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C5 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_15_25_5_30_HV_A4 

VIARULE VIA06_GEN_15_25_10_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C5 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_15_25_10_30_HV_A4 

VIARULE VIA06_GEN_15_25_15_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C5 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_15_25_15_30_HV_A4 

VIARULE VIA06_GEN_15_25_20_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.025 0.015 ;
  LAYER C5 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_15_25_20_30_HV_A4 

VIARULE VIA06_GEN_20_20_0_32_XV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_20_0_32_XV_A4 

VIARULE VIA06_GEN_20_20_2_32_XV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_20_2_32_XV_A4 

VIARULE VIA06_GEN_20_20_5_30_XV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_20_5_30_XV_A4 

VIARULE VIA06_GEN_20_20_10_30_XV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_20_10_30_XV_A4 

VIARULE VIA06_GEN_20_20_15_30_XV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_20_15_30_XV_A4 

VIARULE VIA06_GEN_20_20_20_30_XV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.020 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_20_20_30_XV_A4 

VIARULE VIA06_GEN_20_30_0_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.000 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_30_0_32_HV_A4 

VIARULE VIA06_GEN_20_30_2_32_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.002 0.032 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_30_2_32_HV_A4 

VIARULE VIA06_GEN_20_30_5_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.005 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_30_5_30_HV_A4 

VIARULE VIA06_GEN_20_30_10_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.010 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_30_10_30_HV_A4 

VIARULE VIA06_GEN_20_30_15_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.015 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_30_15_30_HV_A4 

VIARULE VIA06_GEN_20_30_20_30_HV_A4 GENERATE
  LAYER C4 ;
    ENCLOSURE 0.030 0.020 ;
  LAYER C5 ;
    ENCLOSURE 0.020 0.030 ;
  LAYER A4 ;
    RECT -0.022 -0.022 0.022 0.022 ;
    SPACING 0.125 BY 0.134 ;
END  VIA06_GEN_20_30_20_30_HV_A4 

#------------------------------------------------------------
#  YS VIA SECTION 
#------------------------------------------------------------
 VIA VIA07 DEFAULT
 LAYER YS ;
 RECT -0.207 -0.207 0.207 0.207 ;
 LAYER C5 ;
 RECT -0.225 -0.279 0.225 0.279 ;
 LAYER JA ;
 RECT -0.279 -0.225 0.279 0.225 ;
 END VIA07
 
 VIA VIA07_18_72_18_72_VV_YS DEFAULT
 LAYER YS ;
 RECT -0.207 -0.207 0.207 0.207 ;
 LAYER C5 ;
 RECT -0.225 -0.279 0.225 0.279 ;
 LAYER JA ;
 RECT -0.225 -0.279 0.225 0.279 ;
 END VIA07_18_72_18_72_VV_YS
 
 VIA VIA07_18_72_18_72_VH_2CUT_H_YS DEFAULT
 LAYER YS ;
 RECT -0.612 -0.207 -0.198 0.207 ;
 RECT 0.198 -0.207 0.612 0.207 ;
 LAYER C5 ;
 RECT -0.630 -0.279 0.630 0.279 ;
 LAYER JA ;
 RECT -0.684 -0.225 0.684 0.225 ;
 END VIA07_18_72_18_72_VH_2CUT_H_YS
 
 VIA VIA07_18_72_18_72_VH_2CUT_V_YS DEFAULT
 LAYER YS ;
 RECT -0.207 -0.612 0.207 -0.198 ;
 RECT -0.207 0.198 0.207 0.612 ;
 LAYER C5 ;
 RECT -0.225 -0.684 0.225 0.684 ;
 LAYER JA ;
 RECT -0.279 -0.630 0.279 0.630 ;
 END VIA07_18_72_18_72_VH_2CUT_V_YS
 
 VIA VIA07_18_72_18_72_VH_4CUT_YS DEFAULT
 LAYER YS ;
 RECT -0.612 -0.612 -0.198 -0.198 ;
 RECT 0.198 -0.612 0.612 -0.198 ;
 RECT -0.612 0.198 -0.198 0.612 ;
 RECT 0.198 0.198 0.612 0.612 ;
 LAYER C5 ;
 RECT -0.630 -0.684 0.630 0.684 ;
 LAYER JA ;
 RECT -0.684 -0.630 0.684 0.630 ;
 END VIA07_18_72_18_72_VH_4CUT_YS
 
VIARULE VIA07_GEN_18_72_18_72_VH_YS GENERATE
  LAYER C5 ;
    ENCLOSURE 0.018 0.072 ;
  LAYER JA ;
    ENCLOSURE 0.072 0.018 ;
  LAYER YS ;
    RECT -0.207 -0.207 0.207 0.207 ;
    SPACING 0.810 BY 0.810 ;
END  VIA07_GEN_18_72_18_72_VH_YS 

#------------------------------------------------------------
#  JV VIA SECTION 
#------------------------------------------------------------
 VIA VIA08 DEFAULT
 LAYER JV ;
 RECT -0.600 -0.600 0.600 0.600 ;
 LAYER JA ;
 RECT -0.900 -1.200 0.900 1.200 ;
 LAYER QA ;
 RECT -1.200 -0.900 1.200 0.900 ;
 END VIA08
 
VIARULE VIA08_GEN_600_300_600_300_HH_JV GENERATE
  LAYER JA ;
    ENCLOSURE 0.300 0.600 ;
  LAYER QA ;
    ENCLOSURE 0.300 0.600 ;
  LAYER JV ;
    RECT -0.600 -0.600 0.600 0.600 ;
    SPACING 1.200 BY 1.200 ;
END  VIA08_GEN_600_300_600_300_HH_JV 

VIARULE VIA08_GEN_600_300_600_300_HV_JV GENERATE
  LAYER JA ;
    ENCLOSURE 0.300 0.600 ;
  LAYER QA ;
    ENCLOSURE 0.600 0.300 ;
  LAYER JV ;
    RECT -0.600 -0.600 0.600 0.600 ;
    SPACING 1.200 BY 1.200 ;
END  VIA08_GEN_600_300_600_300_HV_JV 

VIARULE VIA08_GEN_600_300_600_300_VH_JV GENERATE
  LAYER JA ;
    ENCLOSURE 0.600 0.300 ;
  LAYER QA ;
    ENCLOSURE 0.300 0.600 ;
  LAYER JV ;
    RECT -0.600 -0.600 0.600 0.600 ;
    SPACING 1.200 BY 1.200 ;
END  VIA08_GEN_600_300_600_300_VH_JV 

VIARULE VIA08_GEN_600_300_600_300_VV_JV GENERATE
  LAYER JA ;
    ENCLOSURE 0.600 0.300 ;
  LAYER QA ;
    ENCLOSURE 0.600 0.300 ;
  LAYER JV ;
    RECT -0.600 -0.600 0.600 0.600 ;
    SPACING 1.200 BY 1.200 ;
END  VIA08_GEN_600_300_600_300_VV_JV 

#------------------------------------------------------------
#  JW VIA SECTION 
#------------------------------------------------------------
 VIA VIA09 DEFAULT
 LAYER JW ;
 RECT -0.600 -0.600 0.600 0.600 ;
 LAYER QA ;
 RECT -1.200 -0.900 1.200 0.900 ;
 LAYER QB ;
 RECT -0.900 -1.200 0.900 1.200 ;
 END VIA09
 
VIARULE VIA09_GEN_600_300_600_300_HH_JW GENERATE
  LAYER QA ;
    ENCLOSURE 0.300 0.600 ;
  LAYER QB ;
    ENCLOSURE 0.300 0.600 ;
  LAYER JW ;
    RECT -0.600 -0.600 0.600 0.600 ;
    SPACING 1.200 BY 1.200 ;
END  VIA09_GEN_600_300_600_300_HH_JW 

VIARULE VIA09_GEN_600_300_600_300_HV_JW GENERATE
  LAYER QA ;
    ENCLOSURE 0.300 0.600 ;
  LAYER QB ;
    ENCLOSURE 0.600 0.300 ;
  LAYER JW ;
    RECT -0.600 -0.600 0.600 0.600 ;
    SPACING 1.200 BY 1.200 ;
END  VIA09_GEN_600_300_600_300_HV_JW 

VIARULE VIA09_GEN_600_300_600_300_VH_JW GENERATE
  LAYER QA ;
    ENCLOSURE 0.600 0.300 ;
  LAYER QB ;
    ENCLOSURE 0.300 0.600 ;
  LAYER JW ;
    RECT -0.600 -0.600 0.600 0.600 ;
    SPACING 1.200 BY 1.200 ;
END  VIA09_GEN_600_300_600_300_VH_JW 

VIARULE VIA09_GEN_600_300_600_300_VV_JW GENERATE
  LAYER QA ;
    ENCLOSURE 0.600 0.300 ;
  LAYER QB ;
    ENCLOSURE 0.600 0.300 ;
  LAYER JW ;
    RECT -0.600 -0.600 0.600 0.600 ;
    SPACING 1.200 BY 1.200 ;
END  VIA09_GEN_600_300_600_300_VV_JW 

#------------------------------------------------------------
#  VV VIA SECTION 
#------------------------------------------------------------
 VIA VIA10 DEFAULT
 LAYER VV ;
 RECT -1.350 -1.350 1.350 1.350 ;
 LAYER QB ;
 RECT -1.800 -1.800 1.800 1.800 ;
 LAYER LB ;
 RECT -1.800 -1.800 1.800 1.800 ;
 END VIA10
 
VIARULE VIA10_GEN_450_450_450_450_XX_VV GENERATE
  LAYER QB ;
    ENCLOSURE 0.450 0.450 ;
  LAYER LB ;
    ENCLOSURE 0.450 0.450 ;
  LAYER VV ;
    RECT -1.350 -1.350 1.350 1.350 ;
    SPACING 4.500 BY 4.500 ;
END  VIA10_GEN_450_450_450_450_XX_VV 


#------------------------------------------------------------------------------
# Special Multi-CUT vias for PG and Bias routing in 6,75 track SNPS IP RFL
#------------------------------------------------------------------------------

VIA VIA01_0_60_0_60_HH_3CUT_H_V1 DEFAULT
LAYER V1 ;
RECT -0.020 -0.020  0.020 0.020 ;
RECT  0.190 -0.020  0.150 0.020 ;
RECT -0.190 -0.020 -0.150 0.020 ;
LAYER M1 ;
RECT -0.250 -0.020 0.250 0.020 ;
LAYER M2 ;
RECT -0.250 -0.020 0.250 0.020 ;
END VIA01_0_60_0_60_HH_3CUT_H_V1

VIA VIA02_0_60_30_60_HH_3CUT_H_AY  DEFAULT
LAYER AY ;
RECT -0.020 -0.020  0.020 0.020 ;
RECT  0.190 -0.020  0.150 0.020 ;
RECT -0.190 -0.020 -0.150 0.020 ;
LAYER M2 ;
RECT -0.250 -0.020 0.250 0.020 ;
LAYER C1 ;
RECT -0.250 -0.050 0.250 0.050 ;
END VIA02_0_60_30_60_HH_3CUT_H_AY

VIA VIA01_0_30_0_30_HH_2CUT_H_V1 DEFAULT
LAYER V1 ;
RECT -0.132 -0.020 -0.092 0.020 ;
RECT  0.092 -0.020  0.132 0.020 ;
LAYER M1 ;
RECT -0.162 -0.020  0.162 0.020 ;
LAYER M2 ;
RECT -0.162 -0.020  0.162 0.020 ;
END VIA01_0_30_0_30_HH_2CUT_H_V1

VIA VIA02_0_30_2_34_HH_2CUT_H_AY DEFAULT
LAYER AY ;
RECT -0.085 -0.020 -0.045 0.020 ;
RECT  0.045 -0.020  0.085 0.020 ;
LAYER M2 ;
RECT -0.115 -0.020 0.115 0.020 ;    
LAYER C1 ;
RECT -0.119 -0.022 0.119 0.022 ;
END VIA02_0_30_2_34_HH_2CUT_H_AY

VIA VIA03_0_41_0_53_HH_2CUT_H_A1 DEFAULT
LAYER A1 ;
RECT -0.085 -0.022 -0.041 0.022 ;
RECT 0.041 -0.022  0.085 0.022 ;
LAYER C1 ;
RECT -0.126 -0.022  0.126 0.022 ;    
LAYER C2 ;
RECT -0.138 -0.022  0.138 0.022 ;
END VIA03_0_41_0_53_HH_2CUT_H_A1

VIA VIA03_BAR_V_0_80_0_80_V_A1 DEFAULT
LAYER A1 ;
RECT -0.022 -0.045 0.022 0.045 ;
LAYER C1 ;
RECT -0.022 -0.125 0.022 0.125 ;
LAYER C2 ;
RECT -0.022 -0.125 0.022 0.125 ;
END VIA03_BAR_V_0_80_0_80_V_A1  

VIA VIA03_32_16_32_16_HH_2CUT_V_A1 DEFAULT
LAYER A1 ;
RECT -0.022 -0.089 0.022 -0.045 ;
RECT -0.022  0.045 0.022  0.089 ;
LAYER C1 ;
RECT -0.054 -0.105 0.054 0.105 ;
LAYER C2 ;
RECT -0.054 -0.105 0.054 0.105 ;
END VIA03_32_16_32_16_HH_2CUT_V_A1

#------------------------------------------------------------------------------

END LIBRARY
