`timescale 1ns/1ps
`define HALF_CLK_CYCLE #10
`define SCAN_DELAY #50

module testbench();

    // Scan chain
    reg phi, phib, scan_i0o1, load, scan_in;
    wire scan_out;

    // Other IO's
    reg clk;
    reg rstn;
    reg reset;
    reg start;
    
    wire clk_div_1k;
    wire [7:0] counter_out;

    // Powers
    supply1 VDD;
    supply1 VDD_TEST;
    supply1 CVDD;
    supply1 DVDD;
    supply0 VSS;

// ==== Extracted from autogenerated testbench by script in tb_scan_chain
   
   // Scan Registers and Initializations
   
`define SCAN_CHAIN_LENGTH 19

   reg [8-1:0] sram_dout;
   reg [8-1:0] sram_dout_read;
   initial sram_dout      = 8'd0;
   initial sram_dout_read = 8'd0;
   reg [1-1:0] en_int;
   reg [1-1:0] en_int_read;
   initial en_int      = 1'd0;
   initial en_int_read = 1'd0;
   reg [1-1:0] en_cnt;
   reg [1-1:0] en_cnt_read;
   initial en_cnt      = 1'd0;
   initial en_cnt_read = 1'd0;
   reg [5-1:0] fc;
   reg [5-1:0] fc_read;
   initial fc      = 5'd0;
   initial fc_read = 5'd0;
   reg [4-1:0] div;
   reg [4-1:0] div_read;
   initial div      = 4'd0;
   initial div_read = 4'd0;
   
   // Scan chain tasks
   
   task load_chip;
      begin
         `SCAN_DELAY load = 1;
         `SCAN_DELAY load = 0;
      end
   endtask

   task load_chain;
      begin
         `SCAN_DELAY scan_i0o1 = 1;
         `SCAN_DELAY phi = 1;
         `SCAN_DELAY phi = 0;
         `SCAN_DELAY phib = 1;
         `SCAN_DELAY phib = 0;
         `SCAN_DELAY scan_i0o1 = 0;
      end
   endtask

   task rotate_chain;
      
      integer i;
      
      reg [`SCAN_CHAIN_LENGTH-1:0] data_in;
      reg [`SCAN_CHAIN_LENGTH-1:0] data_out;
      
      begin
         data_in[7:0] = sram_dout;
         data_in[8:8] = en_int;
         data_in[9:9] = en_cnt;
         data_in[14:10] = fc;
         data_in[18:15] = div;

         for (i = 0; i < `SCAN_CHAIN_LENGTH; i=i+1) begin
            scan_in = data_in[`SCAN_CHAIN_LENGTH-1];
            data_out     = {data_out[`SCAN_CHAIN_LENGTH-2:0], scan_out};
            `SCAN_DELAY phi = 1;
            `SCAN_DELAY phi = 0;
            `SCAN_DELAY phib = 1;
            `SCAN_DELAY phib = 0;
            `SCAN_DELAY data_in = data_in << 1;
         end

         sram_dout_read = data_out[7:0];
         en_int_read = data_out[8:8];
         en_cnt_read = data_out[9:9];
         fc_read = data_out[14:10];
         div_read = data_out[18:15];
      end
      
   endtask

// ====

    chip chip_inst (
        .VDD(VDD), 
	    .VDD_TEST(VDD_TEST), 
	    .CVDD(CVDD), 
	    .DVDD(DVDD), 
	    .VSS(VSS), 
	    
        .BD_to_PAD_phi(phi), 
	    .BD_to_PAD_phib(phib), 
	    .BD_to_PAD_scan_i0o1(scan_i0o1), 
	    .BD_to_PAD_load(load), 
	    .BD_to_PAD_scan_in(scan_in), 
	    .PAD_to_BD_scan_out(scan_out),

	    .BD_to_PAD_clk_ext(clk), 
	    .BD_to_PAD_rstn(rstn), 
	    .BD_to_PAD_reset(reset), 
	    .BD_to_PAD_start(start), 
	    .PAD_to_BD_clk_div_1k(clk_div_1k), 
	    .PAD_to_BD_counter_out(counter_out)
    );

    always begin
        `HALF_CLK_CYCLE clk = ~clk;
    end

    initial begin
        
        //$dumpfile("./vcd_files/chip.vcd");
        //$dumpvars(0, testbench.chip_inst);
        
        // Intialize
        phi=0;
	    phib=0;
	    scan_i0o1=0;
	    load=0;
	    scan_in=0;
        
        clk = 1'b0;
        rstn = 1'b0;
        reset = 1'b0;
        start = 1'b0;
       
        // Scan in initialized value
        rotate_chain();
        load_chip();
        
        // Set values to scan in 
        en_int = 1'b1;
        en_cnt = 1'b1;
        fc = 10;
        div = 3;
       
        // Scan in
        rotate_chain();
        load_chip();

        // global reset
        @(negedge clk);
        rstn = 1'b1;
        @(negedge clk);
        rstn = 1'b0;
        @(negedge clk);
        rstn = 1'b1;
        @(posedge clk);
        @(posedge clk);
    
        // start counting
        @(negedge clk);
        start = 1'b1;
        repeat(500) @(posedge clk);

        // reset
        @(negedge clk);
        start = 1'b0; 
        @(negedge clk);
        reset = 1'b1;
        @(negedge clk);
        @(negedge clk);
        @(negedge clk);
        reset = 1'b0;
        @(negedge clk);
        @(negedge clk);
        @(negedge clk);
        start = 1'b1; 
        repeat(500) @(posedge clk);
       
        // Scan out
        load_chain();
        rotate_chain();
        repeat(500) @(posedge clk);

        //$dumpall;
        //$dumpflush;
        
        $finish;
    end

endmodule
