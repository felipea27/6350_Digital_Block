

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO TOP 
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.00416 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.000208 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.020424 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.000772 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 2.03068 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.09201 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.33792 LAYER C2 ; 
    ANTENNAMAXAREACAR 31.189 LAYER C2 ;
    ANTENNAMAXSIDEAREACAR 1.42437 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 0.005896 LAYER A2 ;
    ANTENNAMAXCUTCAR 1.20182 LAYER A2 ;
    ANTENNAPARTIALMETALAREA 0.845156 LAYER C3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.038068 LAYER C3 ;
    ANTENNAGATEAREA 1.536 LAYER C3 ; 
    ANTENNAMAXAREACAR 41.1563 LAYER C3 ;
    ANTENNAMAXSIDEAREACAR 2.00489 LAYER C3 ;
    ANTENNAPARTIALCUTAREA 0.003872 LAYER A3 ;
    ANTENNAMAXCUTCAR 1.50486 LAYER A3 ;
    ANTENNAPARTIALMETALAREA 0.064944 LAYER C4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003128 LAYER C4 ;
    ANTENNAGATEAREA 1.7664 LAYER C4 ; 
    ANTENNAMAXAREACAR 41.1931 LAYER C4 ;
    ANTENNAMAXSIDEAREACAR 2.00666 LAYER C4 ;
    ANTENNAMAXCUTCAR 1.50486 LAYER A4 ;
  END clk
  PIN rfin 
    ANTENNAPARTIALMETALAREA 0.283976 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.012996 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.006 LAYER C1 ; 
    ANTENNAMAXAREACAR 50.1227 LAYER C1 ;
    ANTENNAMAXSIDEAREACAR 2.296 LAYER C1 ;
    ANTENNAMAXCUTCAR 0.266667 LAYER A1 ;
  END rfin
  PIN rst 
    ANTENNAPARTIALMETALAREA 0.03216 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001608 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0016 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.023364 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00115 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.001936 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.191356 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008874 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 0.005896 LAYER A2 ;
    ANTENNAPARTIALMETALAREA 0.545188 LAYER C3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.024756 LAYER C3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01968 LAYER C3 ; 
    ANTENNAMAXAREACAR 74.2021 LAYER C3 ;
    ANTENNAMAXSIDEAREACAR 3.35246 LAYER C3 ;
    ANTENNAMAXCUTCAR 1.44792 LAYER A3 ;
  END rst
  PIN MOSI 
    ANTENNAPARTIALMETALAREA 0.02216 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.000988 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.661804 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03017 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.144436 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.006452 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.006 LAYER C2 ; 
    ANTENNAMAXAREACAR 33.2847 LAYER C2 ;
    ANTENNAMAXSIDEAREACAR 1.46967 LAYER C2 ;
    ANTENNAMAXCUTCAR 1.19333 LAYER A2 ;
  END MOSI
  PIN CS 
    ANTENNAPARTIALMETALAREA 0.01496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.000628 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.374924 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01713 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.162944 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007092 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.006 LAYER C2 ; 
    ANTENNAMAXAREACAR 38.718 LAYER C2 ;
    ANTENNAMAXSIDEAREACAR 1.72633 LAYER C2 ;
    ANTENNAMAXCUTCAR 1.19333 LAYER A2 ;
  END CS
  PIN SCK 
    ANTENNAPARTIALMETALAREA 0.03296 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001528 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.687324 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03133 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.170864 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007452 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.006 LAYER C2 ; 
    ANTENNAMAXAREACAR 38.0513 LAYER C2 ;
    ANTENNAMAXSIDEAREACAR 1.69067 LAYER C2 ;
    ANTENNAMAXCUTCAR 1.19333 LAYER A2 ;
  END SCK
  PIN TX_BY 
    ANTENNAPARTIALMETALAREA 0.00336 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.000168 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0016 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.277244 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01269 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.001936 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.190872 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008764 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.006 LAYER C2 ; 
    ANTENNAMAXAREACAR 37.4193 LAYER C2 ;
    ANTENNAMAXSIDEAREACAR 1.73633 LAYER C2 ;
    ANTENNAMAXCUTCAR 0.589333 LAYER A2 ;
  END TX_BY
  PIN RX 
    ANTENNAPARTIALMETALAREA 0.02936 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001348 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.339284 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01551 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.139184 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.006012 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.006 LAYER C2 ; 
    ANTENNAMAXAREACAR 80.7713 LAYER C2 ;
    ANTENNAMAXSIDEAREACAR 3.636 LAYER C2 ;
    ANTENNAMAXCUTCAR 1.19333 LAYER A2 ;
  END RX
  PIN pkt_rec 
    ANTENNAPARTIALMETALAREA 0.03656 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001708 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.029524 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00143 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.3845 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.017364 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 0.001936 LAYER A2 ;
    ANTENNAPARTIALMETALAREA 0.011 LAYER C3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.000588 LAYER C3 ;
    ANTENNAPARTIALCUTAREA 0.001936 LAYER A3 ;
    ANTENNAPARTIALMETALAREA 0.349272 LAYER C4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015964 LAYER C4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00672 LAYER C4 ; 
    ANTENNAMAXAREACAR 149.559 LAYER C4 ;
    ANTENNAMAXSIDEAREACAR 6.85536 LAYER C4 ;
    ANTENNAMAXCUTCAR 1.34048 LAYER A4 ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNAGATEAREA 0.01846 LAYER C4 ; 
    ANTENNAMAXAREACAR 65.896 LAYER C4 ;
    ANTENNAMAXSIDEAREACAR 2.96121 LAYER C4 ;
    ANTENNAMAXCUTCAR 0.880607 LAYER A4 ;
  END pkt_rec
  PIN MISO 
    ANTENNAPARTIALMETALAREA 0.01856 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.000808 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.499472 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02259 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.172156 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007712 LAYER C2 ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNAGATEAREA 0.01846 LAYER C2 ; 
    ANTENNAMAXAREACAR 12.9599 LAYER C2 ;
    ANTENNAMAXSIDEAREACAR 0.560888 LAYER C2 ;
    ANTENNAMAXCUTCAR 0.561213 LAYER A2 ;
  END MISO
  PIN TX_OUT 
    ANTENNAPARTIALMETALAREA 0.02496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001248 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0016 LAYER AY ;
    ANTENNAPARTIALMETALAREA 0.021604 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00107 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.001936 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.175032 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008044 LAYER C2 ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNAGATEAREA 0.01846 LAYER C2 ; 
    ANTENNAMAXAREACAR 11.7677 LAYER C2 ;
    ANTENNAMAXSIDEAREACAR 0.513109 LAYER C2 ;
    ANTENNAMAXCUTCAR 0.451571 LAYER A2 ;
  END TX_OUT
  PIN sh_en 
    ANTENNAPARTIALMETALAREA 0.488032 LAYER C1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.021982 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALMETALAREA 0.025636 LAYER C2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001052 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAPARTIALMETALAREA 0.70834 LAYER C3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.032172 LAYER C3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02628 LAYER C3 ; 
    ANTENNAMAXAREACAR 71.0829 LAYER C3 ;
    ANTENNAMAXSIDEAREACAR 3.26205 LAYER C3 ;
    ANTENNAMAXCUTCAR 1.65278 LAYER A3 ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNAGATEAREA 0.00882 LAYER C3 ; 
    ANTENNAMAXAREACAR 111.17 LAYER C3 ;
    ANTENNAMAXSIDEAREACAR 5.00839 LAYER C3 ;
    ANTENNAMAXCUTCAR 1.85029 LAYER A3 ;
  END sh_en
END TOP

END LIBRARY
